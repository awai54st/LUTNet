`timescale 1 ns / 1 ps

module LUTARRAY_32u_1u_s (
        in_V,
        in_1_V,
        in_2_V,
        in_3_V,
        weight_0_V_read,
        ap_return);



input  [63:0] in_V;
input  [63:0] in_1_V;
input  [63:0] in_2_V;
input  [63:0] in_3_V;
input  [63:0] weight_0_V_read;
output  [63:0] ap_return;
wire tmp_0_0;
assign tmp_0_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_V_read[0]);
wire tmp_0_1;
assign tmp_0_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_V_read[1]);
wire tmp_0_2;
assign tmp_0_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_V_read[2]);
wire tmp_0_3;
assign tmp_0_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_V_read[3]);
wire tmp_0_4;
assign tmp_0_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_V_read[4]);
wire tmp_0_5;
assign tmp_0_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_V_read[5]);
wire tmp_0_6;
assign tmp_0_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_V_read[6]);
wire tmp_0_7;
assign tmp_0_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_V_read[7]);
wire tmp_0_8;
assign tmp_0_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_V_read[8]);
wire tmp_0_9;
assign tmp_0_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_V_read[9]);
wire tmp_0_10;
assign tmp_0_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_V_read[10]);
wire tmp_0_11;
assign tmp_0_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_V_read[11]);
wire tmp_0_12;
assign tmp_0_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_V_read[12]);
wire tmp_0_13;
assign tmp_0_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_V_read[13]);
wire tmp_0_14;
assign tmp_0_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_V_read[14]);
wire tmp_0_15;
assign tmp_0_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_V_read[15]);
wire tmp_0_16;
assign tmp_0_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_V_read[16]);
wire tmp_0_17;
assign tmp_0_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_V_read[17]);
wire tmp_0_18;
assign tmp_0_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_V_read[18]);
wire tmp_0_19;
assign tmp_0_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_V_read[19]);
wire tmp_0_20;
assign tmp_0_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_V_read[20]);
wire tmp_0_21;
assign tmp_0_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_V_read[21]);
wire tmp_0_22;
assign tmp_0_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_V_read[22]);
wire tmp_0_23;
assign tmp_0_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_V_read[23]);
wire tmp_0_24;
assign tmp_0_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_V_read[24]);
wire tmp_0_25;
assign tmp_0_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_V_read[25]);
wire tmp_0_26;
assign tmp_0_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_V_read[26]);
wire tmp_0_27;
assign tmp_0_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_V_read[27]);
wire tmp_0_28;
assign tmp_0_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_V_read[28]);
wire tmp_0_29;
assign tmp_0_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_V_read[29]);
wire tmp_0_30;
assign tmp_0_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_V_read[30]);
wire tmp_0_31;
assign tmp_0_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_V_read[31]);
wire tmp_0_32;
assign tmp_0_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_V_read[32]);
wire tmp_0_33;
assign tmp_0_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_V_read[33]);
wire tmp_0_34;
assign tmp_0_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_V_read[34]);
wire tmp_0_35;
assign tmp_0_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_V_read[35]);
wire tmp_0_36;
assign tmp_0_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_V_read[36]);
wire tmp_0_37;
assign tmp_0_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_V_read[37]);
wire tmp_0_38;
assign tmp_0_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_V_read[38]);
wire tmp_0_39;
assign tmp_0_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_V_read[39]);
wire tmp_0_40;
assign tmp_0_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_V_read[40]);
wire tmp_0_41;
assign tmp_0_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_V_read[41]);
wire tmp_0_42;
assign tmp_0_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_V_read[42]);
wire tmp_0_43;
assign tmp_0_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_V_read[43]);
wire tmp_0_44;
assign tmp_0_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_V_read[44]);
wire tmp_0_45;
assign tmp_0_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_V_read[45]);
wire tmp_0_46;
assign tmp_0_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_V_read[46]);
wire tmp_0_47;
assign tmp_0_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_V_read[47]);
wire tmp_0_48;
assign tmp_0_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_V_read[48]);
wire tmp_0_49;
assign tmp_0_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_V_read[49]);
wire tmp_0_50;
assign tmp_0_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_V_read[50]);
wire tmp_0_51;
assign tmp_0_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_V_read[51]);
wire tmp_0_52;
assign tmp_0_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_V_read[52]);
wire tmp_0_53;
assign tmp_0_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_V_read[53]);
wire tmp_0_54;
assign tmp_0_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_V_read[54]);
wire tmp_0_55;
assign tmp_0_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_V_read[55]);
wire tmp_0_56;
assign tmp_0_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_V_read[56]);
wire tmp_0_57;
assign tmp_0_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_V_read[57]);
wire tmp_0_58;
assign tmp_0_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_V_read[58]);
wire tmp_0_59;
assign tmp_0_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_V_read[59]);
wire tmp_0_60;
assign tmp_0_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_V_read[60]);
wire tmp_0_61;
assign tmp_0_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_V_read[61]);
wire tmp_0_62;
assign tmp_0_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_V_read[62]);
wire tmp_0_63;
assign tmp_0_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_V_read[63]);
assign ap_return = {tmp_0_0,tmp_0_1,tmp_0_2,tmp_0_3,tmp_0_4,tmp_0_5,tmp_0_6,tmp_0_7,tmp_0_8,tmp_0_9,tmp_0_10,tmp_0_11,tmp_0_12,tmp_0_13,tmp_0_14,tmp_0_15,tmp_0_16,tmp_0_17,tmp_0_18,tmp_0_19,tmp_0_20,tmp_0_21,tmp_0_22,tmp_0_23,tmp_0_24,tmp_0_25,tmp_0_26,tmp_0_27,tmp_0_28,tmp_0_29,tmp_0_30,tmp_0_31,tmp_0_32,tmp_0_33,tmp_0_34,tmp_0_35,tmp_0_36,tmp_0_37,tmp_0_38,tmp_0_39,tmp_0_40,tmp_0_41,tmp_0_42,tmp_0_43,tmp_0_44,tmp_0_45,tmp_0_46,tmp_0_47,tmp_0_48,tmp_0_49,tmp_0_50,tmp_0_51,tmp_0_52,tmp_0_53,tmp_0_54,tmp_0_55,tmp_0_56,tmp_0_57,tmp_0_58,tmp_0_59,tmp_0_60,tmp_0_61,tmp_0_62,tmp_0_63};
endmodule