`timescale 1 ns / 1 ps

module LUTARRAY_1 (
        in_V,
        in_1_V,
        in_2_V,
        in_3_V,
        weight_0_0_V_read,
        weight_0_1_V_read,
        weight_0_2_V_read,
        weight_0_3_V_read,
        weight_0_4_V_read,
        weight_0_5_V_read,
        weight_0_6_V_read,
        weight_0_7_V_read,
        weight_0_8_V_read,
        weight_0_9_V_read,
        weight_0_10_V_read,
        weight_0_11_V_read,
        weight_0_12_V_read,
        weight_0_13_V_read,
        weight_0_14_V_read,
        weight_0_15_V_read,
        weight_0_16_V_read,
        weight_0_17_V_read,
        weight_0_18_V_read,
        weight_0_19_V_read,
        weight_0_20_V_read,
        weight_0_21_V_read,
        weight_0_22_V_read,
        weight_0_23_V_read,
        weight_0_24_V_read,
        weight_0_25_V_read,
        weight_0_26_V_read,
        weight_0_27_V_read,
        weight_0_28_V_read,
        weight_0_29_V_read,
        weight_0_30_V_read,
        weight_0_31_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31);



input  [31:0] in_V;
input  [31:0] in_1_V;
input  [31:0] in_2_V;
input  [31:0] in_3_V;
input  [31:0] weight_0_0_V_read;
input  [31:0] weight_0_1_V_read;
input  [31:0] weight_0_2_V_read;
input  [31:0] weight_0_3_V_read;
input  [31:0] weight_0_4_V_read;
input  [31:0] weight_0_5_V_read;
input  [31:0] weight_0_6_V_read;
input  [31:0] weight_0_7_V_read;
input  [31:0] weight_0_8_V_read;
input  [31:0] weight_0_9_V_read;
input  [31:0] weight_0_10_V_read;
input  [31:0] weight_0_11_V_read;
input  [31:0] weight_0_12_V_read;
input  [31:0] weight_0_13_V_read;
input  [31:0] weight_0_14_V_read;
input  [31:0] weight_0_15_V_read;
input  [31:0] weight_0_16_V_read;
input  [31:0] weight_0_17_V_read;
input  [31:0] weight_0_18_V_read;
input  [31:0] weight_0_19_V_read;
input  [31:0] weight_0_20_V_read;
input  [31:0] weight_0_21_V_read;
input  [31:0] weight_0_22_V_read;
input  [31:0] weight_0_23_V_read;
input  [31:0] weight_0_24_V_read;
input  [31:0] weight_0_25_V_read;
input  [31:0] weight_0_26_V_read;
input  [31:0] weight_0_27_V_read;
input  [31:0] weight_0_28_V_read;
input  [31:0] weight_0_29_V_read;
input  [31:0] weight_0_30_V_read;
input  [31:0] weight_0_31_V_read;
output  [31:0] ap_return_0;
output  [31:0] ap_return_1;
output  [31:0] ap_return_2;
output  [31:0] ap_return_3;
output  [31:0] ap_return_4;
output  [31:0] ap_return_5;
output  [31:0] ap_return_6;
output  [31:0] ap_return_7;
output  [31:0] ap_return_8;
output  [31:0] ap_return_9;
output  [31:0] ap_return_10;
output  [31:0] ap_return_11;
output  [31:0] ap_return_12;
output  [31:0] ap_return_13;
output  [31:0] ap_return_14;
output  [31:0] ap_return_15;
output  [31:0] ap_return_16;
output  [31:0] ap_return_17;
output  [31:0] ap_return_18;
output  [31:0] ap_return_19;
output  [31:0] ap_return_20;
output  [31:0] ap_return_21;
output  [31:0] ap_return_22;
output  [31:0] ap_return_23;
output  [31:0] ap_return_24;
output  [31:0] ap_return_25;
output  [31:0] ap_return_26;
output  [31:0] ap_return_27;
output  [31:0] ap_return_28;
output  [31:0] ap_return_29;
output  [31:0] ap_return_30;
output  [31:0] ap_return_31;
wire tmp_0_0;
assign tmp_0_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]);
wire tmp_0_1;
assign tmp_0_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]);
wire tmp_0_2;
assign tmp_0_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]);
wire tmp_0_3;
assign tmp_0_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]);
wire tmp_0_4;
assign tmp_0_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]);
wire tmp_0_5;
assign tmp_0_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]);
wire tmp_0_6;
assign tmp_0_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]);
wire tmp_0_7;
assign tmp_0_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]);
wire tmp_0_8;
assign tmp_0_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]);
wire tmp_0_9;
assign tmp_0_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]);
wire tmp_0_10;
assign tmp_0_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]);
wire tmp_0_11;
assign tmp_0_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]);
wire tmp_0_14;
assign tmp_0_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]);
wire tmp_0_15;
assign tmp_0_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]);
wire tmp_0_16;
assign tmp_0_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]);
wire tmp_0_17;
assign tmp_0_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]);
wire tmp_0_18;
assign tmp_0_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]);
wire tmp_0_19;
assign tmp_0_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]);
wire tmp_0_20;
assign tmp_0_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]);
wire tmp_0_21;
assign tmp_0_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]);
wire tmp_0_22;
assign tmp_0_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]);
wire tmp_0_23;
assign tmp_0_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]);
wire tmp_0_24;
assign tmp_0_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]);
wire tmp_0_25;
assign tmp_0_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]);
wire tmp_0_26;
assign tmp_0_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]);
wire tmp_0_27;
assign tmp_0_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]);
wire tmp_0_28;
assign tmp_0_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]);
wire tmp_0_29;
assign tmp_0_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]);
wire tmp_0_30;
assign tmp_0_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]);
wire tmp_0_31;
assign tmp_0_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]);
assign ap_return_0 = {tmp_0_0,tmp_0_1,tmp_0_2,tmp_0_3,tmp_0_4,tmp_0_5,tmp_0_6,tmp_0_7,tmp_0_8,tmp_0_9,tmp_0_10,tmp_0_11,1'b0,1'b0,tmp_0_14,tmp_0_15,tmp_0_16,tmp_0_17,tmp_0_18,tmp_0_19,tmp_0_20,tmp_0_21,tmp_0_22,tmp_0_23,tmp_0_24,tmp_0_25,tmp_0_26,tmp_0_27,tmp_0_28,tmp_0_29,tmp_0_30,tmp_0_31};
wire tmp_1_0;
assign tmp_1_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]);
wire tmp_1_1;
assign tmp_1_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]);
wire tmp_1_2;
assign tmp_1_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]);
wire tmp_1_3;
assign tmp_1_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]);
wire tmp_1_4;
assign tmp_1_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]);
wire tmp_1_5;
assign tmp_1_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]);
wire tmp_1_6;
assign tmp_1_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]);
wire tmp_1_7;
assign tmp_1_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]);
wire tmp_1_9;
assign tmp_1_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]);
wire tmp_1_10;
assign tmp_1_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]);
wire tmp_1_11;
assign tmp_1_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]);
wire tmp_1_12;
assign tmp_1_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]);
wire tmp_1_13;
assign tmp_1_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]);
wire tmp_1_14;
assign tmp_1_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]);
wire tmp_1_15;
assign tmp_1_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]);
wire tmp_1_16;
assign tmp_1_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]);
wire tmp_1_17;
assign tmp_1_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]);
wire tmp_1_18;
assign tmp_1_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]);
wire tmp_1_19;
assign tmp_1_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]);
wire tmp_1_21;
assign tmp_1_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]);
wire tmp_1_23;
assign tmp_1_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]);
wire tmp_1_24;
assign tmp_1_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]);
wire tmp_1_25;
assign tmp_1_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]);
wire tmp_1_26;
assign tmp_1_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]);
wire tmp_1_27;
assign tmp_1_27 = (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]);
wire tmp_1_28;
assign tmp_1_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]);
wire tmp_1_29;
assign tmp_1_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]);
assign ap_return_1 = {tmp_1_0,tmp_1_1,tmp_1_2,tmp_1_3,tmp_1_4,tmp_1_5,tmp_1_6,tmp_1_7,1'b0,tmp_1_9,tmp_1_10,tmp_1_11,tmp_1_12,tmp_1_13,tmp_1_14,tmp_1_15,tmp_1_16,tmp_1_17,tmp_1_18,tmp_1_19,1'b0,tmp_1_21,1'b0,tmp_1_23,tmp_1_24,tmp_1_25,tmp_1_26,tmp_1_27,tmp_1_28,tmp_1_29,1'b0,1'b0};
wire tmp_2_0;
assign tmp_2_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]);
wire tmp_2_1;
assign tmp_2_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]);
wire tmp_2_2;
assign tmp_2_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]);
wire tmp_2_3;
assign tmp_2_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]);
wire tmp_2_4;
assign tmp_2_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]);
wire tmp_2_5;
assign tmp_2_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]);
wire tmp_2_6;
assign tmp_2_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]);
wire tmp_2_7;
assign tmp_2_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]);
wire tmp_2_10;
assign tmp_2_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]);
wire tmp_2_11;
assign tmp_2_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]);
wire tmp_2_12;
assign tmp_2_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]);
wire tmp_2_13;
assign tmp_2_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]);
wire tmp_2_14;
assign tmp_2_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]);
wire tmp_2_15;
assign tmp_2_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]);
wire tmp_2_16;
assign tmp_2_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]);
wire tmp_2_18;
assign tmp_2_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]);
wire tmp_2_19;
assign tmp_2_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]);
wire tmp_2_20;
assign tmp_2_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]);
wire tmp_2_21;
assign tmp_2_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]);
wire tmp_2_22;
assign tmp_2_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]);
wire tmp_2_23;
assign tmp_2_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]);
wire tmp_2_24;
assign tmp_2_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]);
wire tmp_2_25;
assign tmp_2_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]);
wire tmp_2_26;
assign tmp_2_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]);
wire tmp_2_27;
assign tmp_2_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]);
wire tmp_2_28;
assign tmp_2_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]);
wire tmp_2_29;
assign tmp_2_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]);
wire tmp_2_30;
assign tmp_2_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]);
wire tmp_2_31;
assign tmp_2_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]);
assign ap_return_2 = {tmp_2_0,tmp_2_1,tmp_2_2,tmp_2_3,tmp_2_4,tmp_2_5,tmp_2_6,tmp_2_7,1'b0,1'b0,tmp_2_10,tmp_2_11,tmp_2_12,tmp_2_13,tmp_2_14,tmp_2_15,tmp_2_16,1'b0,tmp_2_18,tmp_2_19,tmp_2_20,tmp_2_21,tmp_2_22,tmp_2_23,tmp_2_24,tmp_2_25,tmp_2_26,tmp_2_27,tmp_2_28,tmp_2_29,tmp_2_30,tmp_2_31};
wire tmp_3_0;
assign tmp_3_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]);
wire tmp_3_1;
assign tmp_3_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]);
wire tmp_3_2;
assign tmp_3_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]);
wire tmp_3_3;
assign tmp_3_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]);
wire tmp_3_4;
assign tmp_3_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]);
wire tmp_3_5;
assign tmp_3_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]);
wire tmp_3_6;
assign tmp_3_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]);
wire tmp_3_7;
assign tmp_3_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]);
wire tmp_3_8;
assign tmp_3_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]);
wire tmp_3_9;
assign tmp_3_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]);
wire tmp_3_10;
assign tmp_3_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]);
wire tmp_3_11;
assign tmp_3_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]);
wire tmp_3_12;
assign tmp_3_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]);
wire tmp_3_13;
assign tmp_3_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]);
wire tmp_3_14;
assign tmp_3_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]);
wire tmp_3_15;
assign tmp_3_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]);
wire tmp_3_16;
assign tmp_3_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]);
wire tmp_3_17;
assign tmp_3_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]);
wire tmp_3_18;
assign tmp_3_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]);
wire tmp_3_19;
assign tmp_3_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]);
wire tmp_3_20;
assign tmp_3_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]);
wire tmp_3_21;
assign tmp_3_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]);
wire tmp_3_23;
assign tmp_3_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]);
wire tmp_3_24;
assign tmp_3_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]);
wire tmp_3_25;
assign tmp_3_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]);
wire tmp_3_26;
assign tmp_3_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]);
wire tmp_3_27;
assign tmp_3_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]);
wire tmp_3_28;
assign tmp_3_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]);
wire tmp_3_29;
assign tmp_3_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]);
wire tmp_3_31;
assign tmp_3_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]);
assign ap_return_3 = {tmp_3_0,tmp_3_1,tmp_3_2,tmp_3_3,tmp_3_4,tmp_3_5,tmp_3_6,tmp_3_7,tmp_3_8,tmp_3_9,tmp_3_10,tmp_3_11,tmp_3_12,tmp_3_13,tmp_3_14,tmp_3_15,tmp_3_16,tmp_3_17,tmp_3_18,tmp_3_19,tmp_3_20,tmp_3_21,1'b0,tmp_3_23,tmp_3_24,tmp_3_25,tmp_3_26,tmp_3_27,tmp_3_28,tmp_3_29,1'b0,tmp_3_31};
wire tmp_4_0;
assign tmp_4_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]);
wire tmp_4_1;
assign tmp_4_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]);
wire tmp_4_2;
assign tmp_4_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]);
wire tmp_4_3;
assign tmp_4_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]);
wire tmp_4_4;
assign tmp_4_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]);
wire tmp_4_5;
assign tmp_4_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]);
wire tmp_4_6;
assign tmp_4_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]);
wire tmp_4_7;
assign tmp_4_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]);
wire tmp_4_8;
assign tmp_4_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]);
wire tmp_4_9;
assign tmp_4_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]);
wire tmp_4_10;
assign tmp_4_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]);
wire tmp_4_11;
assign tmp_4_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]);
wire tmp_4_12;
assign tmp_4_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]);
wire tmp_4_13;
assign tmp_4_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]);
wire tmp_4_14;
assign tmp_4_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]);
wire tmp_4_15;
assign tmp_4_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]);
wire tmp_4_16;
assign tmp_4_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]);
wire tmp_4_17;
assign tmp_4_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]);
wire tmp_4_18;
assign tmp_4_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]);
wire tmp_4_19;
assign tmp_4_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]);
wire tmp_4_20;
assign tmp_4_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]);
wire tmp_4_21;
assign tmp_4_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]);
wire tmp_4_22;
assign tmp_4_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]);
wire tmp_4_23;
assign tmp_4_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]);
wire tmp_4_24;
assign tmp_4_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]);
wire tmp_4_25;
assign tmp_4_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]);
wire tmp_4_26;
assign tmp_4_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]);
wire tmp_4_27;
assign tmp_4_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]);
wire tmp_4_28;
assign tmp_4_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]);
wire tmp_4_30;
assign tmp_4_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]);
wire tmp_4_31;
assign tmp_4_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]);
assign ap_return_4 = {tmp_4_0,tmp_4_1,tmp_4_2,tmp_4_3,tmp_4_4,tmp_4_5,tmp_4_6,tmp_4_7,tmp_4_8,tmp_4_9,tmp_4_10,tmp_4_11,tmp_4_12,tmp_4_13,tmp_4_14,tmp_4_15,tmp_4_16,tmp_4_17,tmp_4_18,tmp_4_19,tmp_4_20,tmp_4_21,tmp_4_22,tmp_4_23,tmp_4_24,tmp_4_25,tmp_4_26,tmp_4_27,tmp_4_28,1'b0,tmp_4_30,tmp_4_31};
wire tmp_5_0;
assign tmp_5_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]);
wire tmp_5_1;
assign tmp_5_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]);
wire tmp_5_2;
assign tmp_5_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]);
wire tmp_5_3;
assign tmp_5_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]);
wire tmp_5_4;
assign tmp_5_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]);
wire tmp_5_5;
assign tmp_5_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]);
wire tmp_5_6;
assign tmp_5_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]);
wire tmp_5_8;
assign tmp_5_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]);
wire tmp_5_9;
assign tmp_5_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]);
wire tmp_5_10;
assign tmp_5_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]);
wire tmp_5_11;
assign tmp_5_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]);
wire tmp_5_12;
assign tmp_5_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]);
wire tmp_5_13;
assign tmp_5_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]);
wire tmp_5_15;
assign tmp_5_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]);
wire tmp_5_16;
assign tmp_5_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]);
wire tmp_5_17;
assign tmp_5_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]);
wire tmp_5_18;
assign tmp_5_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]);
wire tmp_5_19;
assign tmp_5_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]);
wire tmp_5_20;
assign tmp_5_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]);
wire tmp_5_21;
assign tmp_5_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]);
wire tmp_5_22;
assign tmp_5_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]);
wire tmp_5_23;
assign tmp_5_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]);
wire tmp_5_24;
assign tmp_5_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]);
wire tmp_5_25;
assign tmp_5_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]);
wire tmp_5_27;
assign tmp_5_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]);
wire tmp_5_28;
assign tmp_5_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]);
wire tmp_5_29;
assign tmp_5_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]);
wire tmp_5_30;
assign tmp_5_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]);
wire tmp_5_31;
assign tmp_5_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]);
assign ap_return_5 = {tmp_5_0,tmp_5_1,tmp_5_2,tmp_5_3,tmp_5_4,tmp_5_5,tmp_5_6,1'b0,tmp_5_8,tmp_5_9,tmp_5_10,tmp_5_11,tmp_5_12,tmp_5_13,1'b0,tmp_5_15,tmp_5_16,tmp_5_17,tmp_5_18,tmp_5_19,tmp_5_20,tmp_5_21,tmp_5_22,tmp_5_23,tmp_5_24,tmp_5_25,1'b0,tmp_5_27,tmp_5_28,tmp_5_29,tmp_5_30,tmp_5_31};
wire tmp_6_0;
assign tmp_6_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]);
wire tmp_6_1;
assign tmp_6_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]);
wire tmp_6_2;
assign tmp_6_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]);
wire tmp_6_3;
assign tmp_6_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]);
wire tmp_6_4;
assign tmp_6_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]);
wire tmp_6_5;
assign tmp_6_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]);
wire tmp_6_6;
assign tmp_6_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]);
wire tmp_6_7;
assign tmp_6_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]);
wire tmp_6_8;
assign tmp_6_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]);
wire tmp_6_9;
assign tmp_6_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]);
wire tmp_6_10;
assign tmp_6_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]);
wire tmp_6_11;
assign tmp_6_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]);
wire tmp_6_12;
assign tmp_6_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]);
wire tmp_6_13;
assign tmp_6_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]);
wire tmp_6_14;
assign tmp_6_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]);
wire tmp_6_15;
assign tmp_6_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]);
wire tmp_6_16;
assign tmp_6_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]);
wire tmp_6_17;
assign tmp_6_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]);
wire tmp_6_18;
assign tmp_6_18 = (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]);
wire tmp_6_19;
assign tmp_6_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]);
wire tmp_6_20;
assign tmp_6_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]);
wire tmp_6_21;
assign tmp_6_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]);
wire tmp_6_22;
assign tmp_6_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]);
wire tmp_6_23;
assign tmp_6_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]);
wire tmp_6_24;
assign tmp_6_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]);
wire tmp_6_26;
assign tmp_6_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]);
wire tmp_6_27;
assign tmp_6_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]);
wire tmp_6_28;
assign tmp_6_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]);
wire tmp_6_29;
assign tmp_6_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]);
wire tmp_6_30;
assign tmp_6_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]);
wire tmp_6_31;
assign tmp_6_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]);
assign ap_return_6 = {tmp_6_0,tmp_6_1,tmp_6_2,tmp_6_3,tmp_6_4,tmp_6_5,tmp_6_6,tmp_6_7,tmp_6_8,tmp_6_9,tmp_6_10,tmp_6_11,tmp_6_12,tmp_6_13,tmp_6_14,tmp_6_15,tmp_6_16,tmp_6_17,tmp_6_18,tmp_6_19,tmp_6_20,tmp_6_21,tmp_6_22,tmp_6_23,tmp_6_24,1'b0,tmp_6_26,tmp_6_27,tmp_6_28,tmp_6_29,tmp_6_30,tmp_6_31};
wire tmp_7_0;
assign tmp_7_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]);
wire tmp_7_1;
assign tmp_7_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]);
wire tmp_7_2;
assign tmp_7_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]);
wire tmp_7_3;
assign tmp_7_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]);
wire tmp_7_4;
assign tmp_7_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]);
wire tmp_7_5;
assign tmp_7_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]);
wire tmp_7_6;
assign tmp_7_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]);
wire tmp_7_7;
assign tmp_7_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]);
wire tmp_7_8;
assign tmp_7_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]);
wire tmp_7_9;
assign tmp_7_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]);
wire tmp_7_10;
assign tmp_7_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]);
wire tmp_7_11;
assign tmp_7_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]);
wire tmp_7_12;
assign tmp_7_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]);
wire tmp_7_13;
assign tmp_7_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]);
wire tmp_7_14;
assign tmp_7_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]);
wire tmp_7_15;
assign tmp_7_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]);
wire tmp_7_16;
assign tmp_7_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]);
wire tmp_7_17;
assign tmp_7_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]);
wire tmp_7_18;
assign tmp_7_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]);
wire tmp_7_19;
assign tmp_7_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]);
wire tmp_7_20;
assign tmp_7_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]);
wire tmp_7_21;
assign tmp_7_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]);
wire tmp_7_22;
assign tmp_7_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]);
wire tmp_7_23;
assign tmp_7_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]);
wire tmp_7_24;
assign tmp_7_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]);
wire tmp_7_25;
assign tmp_7_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]);
wire tmp_7_26;
assign tmp_7_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]);
wire tmp_7_27;
assign tmp_7_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]);
wire tmp_7_28;
assign tmp_7_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]);
wire tmp_7_29;
assign tmp_7_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]);
wire tmp_7_30;
assign tmp_7_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]);
wire tmp_7_31;
assign tmp_7_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]);
assign ap_return_7 = {tmp_7_0,tmp_7_1,tmp_7_2,tmp_7_3,tmp_7_4,tmp_7_5,tmp_7_6,tmp_7_7,tmp_7_8,tmp_7_9,tmp_7_10,tmp_7_11,tmp_7_12,tmp_7_13,tmp_7_14,tmp_7_15,tmp_7_16,tmp_7_17,tmp_7_18,tmp_7_19,tmp_7_20,tmp_7_21,tmp_7_22,tmp_7_23,tmp_7_24,tmp_7_25,tmp_7_26,tmp_7_27,tmp_7_28,tmp_7_29,tmp_7_30,tmp_7_31};
wire tmp_8_0;
assign tmp_8_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]);
wire tmp_8_1;
assign tmp_8_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]);
wire tmp_8_2;
assign tmp_8_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]);
wire tmp_8_3;
assign tmp_8_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]);
wire tmp_8_4;
assign tmp_8_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_8_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_8_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_8_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_8_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_8_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_8_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_8_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_8_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_8_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_8_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_8_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_8_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_8_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_8_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_8_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_8_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_8_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_8_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_8_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_8_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_8_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_8_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_8_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_8_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_8_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_8_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_8_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_8_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_8_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_8_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_8_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_8_V_read[4]);
wire tmp_8_5;
assign tmp_8_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]);
wire tmp_8_6;
assign tmp_8_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]);
wire tmp_8_8;
assign tmp_8_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]);
wire tmp_8_9;
assign tmp_8_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]);
wire tmp_8_10;
assign tmp_8_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]);
wire tmp_8_11;
assign tmp_8_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]);
wire tmp_8_12;
assign tmp_8_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]);
wire tmp_8_13;
assign tmp_8_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]);
wire tmp_8_14;
assign tmp_8_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]);
wire tmp_8_16;
assign tmp_8_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]);
wire tmp_8_17;
assign tmp_8_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]);
wire tmp_8_18;
assign tmp_8_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]);
wire tmp_8_19;
assign tmp_8_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]);
wire tmp_8_20;
assign tmp_8_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]);
wire tmp_8_21;
assign tmp_8_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]);
wire tmp_8_22;
assign tmp_8_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]);
wire tmp_8_23;
assign tmp_8_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]);
wire tmp_8_25;
assign tmp_8_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]);
wire tmp_8_27;
assign tmp_8_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]);
wire tmp_8_28;
assign tmp_8_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]);
wire tmp_8_29;
assign tmp_8_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]);
wire tmp_8_30;
assign tmp_8_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]);
wire tmp_8_31;
assign tmp_8_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]);
assign ap_return_8 = {tmp_8_0,tmp_8_1,tmp_8_2,tmp_8_3,tmp_8_4,tmp_8_5,tmp_8_6,1'b0,tmp_8_8,tmp_8_9,tmp_8_10,tmp_8_11,tmp_8_12,tmp_8_13,tmp_8_14,1'b0,tmp_8_16,tmp_8_17,tmp_8_18,tmp_8_19,tmp_8_20,tmp_8_21,tmp_8_22,tmp_8_23,1'b0,tmp_8_25,1'b0,tmp_8_27,tmp_8_28,tmp_8_29,tmp_8_30,tmp_8_31};
wire tmp_9_0;
assign tmp_9_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]);
wire tmp_9_1;
assign tmp_9_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]);
wire tmp_9_2;
assign tmp_9_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]);
wire tmp_9_3;
assign tmp_9_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]);
wire tmp_9_4;
assign tmp_9_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]);
wire tmp_9_5;
assign tmp_9_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]);
wire tmp_9_6;
assign tmp_9_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_9_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_9_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_9_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_9_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_9_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_9_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_9_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_9_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_9_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_9_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_9_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_9_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_9_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_9_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_9_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_9_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_9_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_9_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_9_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_9_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_9_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_9_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_9_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_9_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_9_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_9_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_9_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_9_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_9_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_9_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_9_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_9_V_read[6]);
wire tmp_9_7;
assign tmp_9_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]);
wire tmp_9_8;
assign tmp_9_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]);
wire tmp_9_9;
assign tmp_9_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]);
wire tmp_9_10;
assign tmp_9_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]);
wire tmp_9_11;
assign tmp_9_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]);
wire tmp_9_12;
assign tmp_9_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]);
wire tmp_9_13;
assign tmp_9_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]);
wire tmp_9_14;
assign tmp_9_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]);
wire tmp_9_15;
assign tmp_9_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]);
wire tmp_9_16;
assign tmp_9_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]);
wire tmp_9_17;
assign tmp_9_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]);
wire tmp_9_18;
assign tmp_9_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]);
wire tmp_9_19;
assign tmp_9_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]);
wire tmp_9_20;
assign tmp_9_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]);
wire tmp_9_22;
assign tmp_9_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]);
wire tmp_9_23;
assign tmp_9_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]);
wire tmp_9_24;
assign tmp_9_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]);
wire tmp_9_25;
assign tmp_9_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]);
wire tmp_9_26;
assign tmp_9_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]);
wire tmp_9_27;
assign tmp_9_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]);
wire tmp_9_28;
assign tmp_9_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]);
wire tmp_9_30;
assign tmp_9_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_9_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_9_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_9_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_9_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_9_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_9_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_9_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_9_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_9_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_9_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_9_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_9_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_9_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_9_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_9_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_9_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_9_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_9_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_9_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_9_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_9_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_9_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_9_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_9_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_9_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_9_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_9_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_9_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_9_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_9_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_9_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_9_V_read[30]);
wire tmp_9_31;
assign tmp_9_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]);
assign ap_return_9 = {tmp_9_0,tmp_9_1,tmp_9_2,tmp_9_3,tmp_9_4,tmp_9_5,tmp_9_6,tmp_9_7,tmp_9_8,tmp_9_9,tmp_9_10,tmp_9_11,tmp_9_12,tmp_9_13,tmp_9_14,tmp_9_15,tmp_9_16,tmp_9_17,tmp_9_18,tmp_9_19,tmp_9_20,1'b0,tmp_9_22,tmp_9_23,tmp_9_24,tmp_9_25,tmp_9_26,tmp_9_27,tmp_9_28,1'b0,tmp_9_30,tmp_9_31};
wire tmp_10_0;
assign tmp_10_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]);
wire tmp_10_1;
assign tmp_10_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]);
wire tmp_10_2;
assign tmp_10_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]);
wire tmp_10_3;
assign tmp_10_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]);
wire tmp_10_4;
assign tmp_10_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]);
wire tmp_10_5;
assign tmp_10_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]);
wire tmp_10_6;
assign tmp_10_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]);
wire tmp_10_7;
assign tmp_10_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]);
wire tmp_10_8;
assign tmp_10_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]);
wire tmp_10_9;
assign tmp_10_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]);
wire tmp_10_10;
assign tmp_10_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]);
wire tmp_10_11;
assign tmp_10_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]);
wire tmp_10_12;
assign tmp_10_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]);
wire tmp_10_13;
assign tmp_10_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]);
wire tmp_10_14;
assign tmp_10_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]);
wire tmp_10_15;
assign tmp_10_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]);
wire tmp_10_16;
assign tmp_10_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]);
wire tmp_10_17;
assign tmp_10_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]);
wire tmp_10_18;
assign tmp_10_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_10_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_10_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_10_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_10_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_10_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_10_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_10_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_10_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_10_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_10_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_10_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_10_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_10_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_10_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_10_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_10_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_10_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_10_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_10_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_10_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_10_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_10_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_10_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_10_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_10_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_10_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_10_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_10_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_10_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_10_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_10_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_10_V_read[18]);
wire tmp_10_19;
assign tmp_10_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]);
wire tmp_10_20;
assign tmp_10_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]);
wire tmp_10_21;
assign tmp_10_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]);
wire tmp_10_22;
assign tmp_10_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]);
wire tmp_10_23;
assign tmp_10_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]);
wire tmp_10_24;
assign tmp_10_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]);
wire tmp_10_25;
assign tmp_10_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]);
wire tmp_10_26;
assign tmp_10_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]);
wire tmp_10_27;
assign tmp_10_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]);
wire tmp_10_28;
assign tmp_10_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]);
wire tmp_10_29;
assign tmp_10_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]);
wire tmp_10_30;
assign tmp_10_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]);
wire tmp_10_31;
assign tmp_10_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]);
assign ap_return_10 = {tmp_10_0,tmp_10_1,tmp_10_2,tmp_10_3,tmp_10_4,tmp_10_5,tmp_10_6,tmp_10_7,tmp_10_8,tmp_10_9,tmp_10_10,tmp_10_11,tmp_10_12,tmp_10_13,tmp_10_14,tmp_10_15,tmp_10_16,tmp_10_17,tmp_10_18,tmp_10_19,tmp_10_20,tmp_10_21,tmp_10_22,tmp_10_23,tmp_10_24,tmp_10_25,tmp_10_26,tmp_10_27,tmp_10_28,tmp_10_29,tmp_10_30,tmp_10_31};
wire tmp_11_0;
assign tmp_11_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]);
wire tmp_11_1;
assign tmp_11_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]);
wire tmp_11_2;
assign tmp_11_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]);
wire tmp_11_3;
assign tmp_11_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]);
wire tmp_11_4;
assign tmp_11_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]);
wire tmp_11_5;
assign tmp_11_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]);
wire tmp_11_6;
assign tmp_11_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]);
wire tmp_11_7;
assign tmp_11_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]);
wire tmp_11_8;
assign tmp_11_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]);
wire tmp_11_9;
assign tmp_11_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]);
wire tmp_11_10;
assign tmp_11_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]);
wire tmp_11_12;
assign tmp_11_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]);
wire tmp_11_13;
assign tmp_11_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]);
wire tmp_11_14;
assign tmp_11_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]);
wire tmp_11_15;
assign tmp_11_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]);
wire tmp_11_16;
assign tmp_11_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]);
wire tmp_11_17;
assign tmp_11_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]);
wire tmp_11_18;
assign tmp_11_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]);
wire tmp_11_19;
assign tmp_11_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]);
wire tmp_11_20;
assign tmp_11_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]);
wire tmp_11_21;
assign tmp_11_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]);
wire tmp_11_22;
assign tmp_11_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]);
wire tmp_11_23;
assign tmp_11_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_11_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_11_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_11_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_11_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_11_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_11_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_11_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_11_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_11_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_11_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_11_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_11_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_11_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_11_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_11_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_11_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_11_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_11_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_11_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_11_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_11_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_11_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_11_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_11_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_11_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_11_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_11_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_11_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_11_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_11_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_11_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_11_V_read[23]);
wire tmp_11_24;
assign tmp_11_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]);
wire tmp_11_25;
assign tmp_11_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_11_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_11_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_11_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_11_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_11_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_11_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_11_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_11_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_11_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_11_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_11_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_11_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_11_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_11_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_11_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_11_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_11_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_11_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_11_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_11_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_11_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_11_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_11_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_11_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_11_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_11_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_11_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_11_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_11_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_11_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_11_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_11_V_read[25]);
wire tmp_11_26;
assign tmp_11_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]);
wire tmp_11_27;
assign tmp_11_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]);
wire tmp_11_28;
assign tmp_11_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]);
wire tmp_11_29;
assign tmp_11_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]);
wire tmp_11_30;
assign tmp_11_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]);
wire tmp_11_31;
assign tmp_11_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]);
assign ap_return_11 = {tmp_11_0,tmp_11_1,tmp_11_2,tmp_11_3,tmp_11_4,tmp_11_5,tmp_11_6,tmp_11_7,tmp_11_8,tmp_11_9,tmp_11_10,1'b0,tmp_11_12,tmp_11_13,tmp_11_14,tmp_11_15,tmp_11_16,tmp_11_17,tmp_11_18,tmp_11_19,tmp_11_20,tmp_11_21,tmp_11_22,tmp_11_23,tmp_11_24,tmp_11_25,tmp_11_26,tmp_11_27,tmp_11_28,tmp_11_29,tmp_11_30,tmp_11_31};
wire tmp_12_0;
assign tmp_12_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]);
wire tmp_12_1;
assign tmp_12_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]);
wire tmp_12_2;
assign tmp_12_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]);
wire tmp_12_3;
assign tmp_12_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]);
wire tmp_12_4;
assign tmp_12_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]);
wire tmp_12_6;
assign tmp_12_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]);
wire tmp_12_7;
assign tmp_12_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]);
wire tmp_12_8;
assign tmp_12_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]);
wire tmp_12_9;
assign tmp_12_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]);
wire tmp_12_10;
assign tmp_12_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]);
wire tmp_12_11;
assign tmp_12_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]);
wire tmp_12_12;
assign tmp_12_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]);
wire tmp_12_13;
assign tmp_12_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]);
wire tmp_12_14;
assign tmp_12_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]);
wire tmp_12_16;
assign tmp_12_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]);
wire tmp_12_17;
assign tmp_12_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]);
wire tmp_12_18;
assign tmp_12_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]);
wire tmp_12_19;
assign tmp_12_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]);
wire tmp_12_21;
assign tmp_12_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]);
wire tmp_12_22;
assign tmp_12_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]);
wire tmp_12_23;
assign tmp_12_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]);
wire tmp_12_24;
assign tmp_12_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]);
wire tmp_12_25;
assign tmp_12_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]);
wire tmp_12_26;
assign tmp_12_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]);
wire tmp_12_27;
assign tmp_12_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]);
wire tmp_12_28;
assign tmp_12_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]);
wire tmp_12_29;
assign tmp_12_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]);
wire tmp_12_30;
assign tmp_12_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]);
wire tmp_12_31;
assign tmp_12_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]);
assign ap_return_12 = {tmp_12_0,tmp_12_1,tmp_12_2,tmp_12_3,tmp_12_4,1'b0,tmp_12_6,tmp_12_7,tmp_12_8,tmp_12_9,tmp_12_10,tmp_12_11,tmp_12_12,tmp_12_13,tmp_12_14,1'b0,tmp_12_16,tmp_12_17,tmp_12_18,tmp_12_19,1'b0,tmp_12_21,tmp_12_22,tmp_12_23,tmp_12_24,tmp_12_25,tmp_12_26,tmp_12_27,tmp_12_28,tmp_12_29,tmp_12_30,tmp_12_31};
wire tmp_13_0;
assign tmp_13_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]);
wire tmp_13_1;
assign tmp_13_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]);
wire tmp_13_2;
assign tmp_13_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]);
wire tmp_13_3;
assign tmp_13_3 = (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]);
wire tmp_13_4;
assign tmp_13_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]);
wire tmp_13_5;
assign tmp_13_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]);
wire tmp_13_6;
assign tmp_13_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_13_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_13_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_13_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_13_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_13_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_13_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_13_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_13_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_13_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_13_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_13_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_13_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_13_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_13_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_13_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_13_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_13_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_13_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_13_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_13_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_13_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_13_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_13_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_13_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_13_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_13_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_13_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_13_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_13_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_13_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_13_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_13_V_read[6]);
wire tmp_13_7;
assign tmp_13_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]);
wire tmp_13_8;
assign tmp_13_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]);
wire tmp_13_9;
assign tmp_13_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]);
wire tmp_13_10;
assign tmp_13_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]);
wire tmp_13_11;
assign tmp_13_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]);
wire tmp_13_12;
assign tmp_13_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]);
wire tmp_13_13;
assign tmp_13_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]);
wire tmp_13_14;
assign tmp_13_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]);
wire tmp_13_15;
assign tmp_13_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]);
wire tmp_13_16;
assign tmp_13_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]);
wire tmp_13_17;
assign tmp_13_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]);
wire tmp_13_18;
assign tmp_13_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]);
wire tmp_13_19;
assign tmp_13_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]);
wire tmp_13_20;
assign tmp_13_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]);
wire tmp_13_21;
assign tmp_13_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]);
wire tmp_13_22;
assign tmp_13_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]);
wire tmp_13_23;
assign tmp_13_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]);
wire tmp_13_24;
assign tmp_13_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]);
wire tmp_13_25;
assign tmp_13_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]);
wire tmp_13_26;
assign tmp_13_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]);
wire tmp_13_27;
assign tmp_13_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]);
wire tmp_13_28;
assign tmp_13_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]);
wire tmp_13_29;
assign tmp_13_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]);
wire tmp_13_31;
assign tmp_13_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]);
assign ap_return_13 = {tmp_13_0,tmp_13_1,tmp_13_2,tmp_13_3,tmp_13_4,tmp_13_5,tmp_13_6,tmp_13_7,tmp_13_8,tmp_13_9,tmp_13_10,tmp_13_11,tmp_13_12,tmp_13_13,tmp_13_14,tmp_13_15,tmp_13_16,tmp_13_17,tmp_13_18,tmp_13_19,tmp_13_20,tmp_13_21,tmp_13_22,tmp_13_23,tmp_13_24,tmp_13_25,tmp_13_26,tmp_13_27,tmp_13_28,tmp_13_29,1'b0,tmp_13_31};
wire tmp_14_0;
assign tmp_14_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]);
wire tmp_14_1;
assign tmp_14_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]);
wire tmp_14_2;
assign tmp_14_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]);
wire tmp_14_3;
assign tmp_14_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]);
wire tmp_14_4;
assign tmp_14_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]);
wire tmp_14_6;
assign tmp_14_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]);
wire tmp_14_7;
assign tmp_14_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]);
wire tmp_14_8;
assign tmp_14_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]);
wire tmp_14_9;
assign tmp_14_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]);
wire tmp_14_10;
assign tmp_14_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]);
wire tmp_14_11;
assign tmp_14_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]);
wire tmp_14_12;
assign tmp_14_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]);
wire tmp_14_13;
assign tmp_14_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]);
wire tmp_14_14;
assign tmp_14_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_14_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_14_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_14_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_14_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_14_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_14_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_14_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_14_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_14_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_14_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_14_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_14_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_14_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_14_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_14_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_14_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_14_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_14_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_14_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_14_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_14_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_14_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_14_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_14_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_14_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_14_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_14_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_14_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_14_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_14_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_14_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_14_V_read[14]);
wire tmp_14_16;
assign tmp_14_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]);
wire tmp_14_17;
assign tmp_14_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]);
wire tmp_14_18;
assign tmp_14_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]);
wire tmp_14_19;
assign tmp_14_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]);
wire tmp_14_20;
assign tmp_14_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]);
wire tmp_14_21;
assign tmp_14_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]);
wire tmp_14_22;
assign tmp_14_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]);
wire tmp_14_23;
assign tmp_14_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]);
wire tmp_14_24;
assign tmp_14_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]);
wire tmp_14_25;
assign tmp_14_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]);
wire tmp_14_26;
assign tmp_14_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]);
wire tmp_14_27;
assign tmp_14_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]);
wire tmp_14_28;
assign tmp_14_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]);
wire tmp_14_29;
assign tmp_14_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]);
wire tmp_14_30;
assign tmp_14_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]);
wire tmp_14_31;
assign tmp_14_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_14_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_14_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_14_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_14_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_14_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_14_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_14_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_14_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_14_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_14_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_14_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_14_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_14_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_14_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_14_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_14_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_14_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_14_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_14_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_14_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_14_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_14_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_14_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_14_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_14_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_14_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_14_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_14_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_14_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_14_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_14_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_14_V_read[31]);
assign ap_return_14 = {tmp_14_0,tmp_14_1,tmp_14_2,tmp_14_3,tmp_14_4,1'b0,tmp_14_6,tmp_14_7,tmp_14_8,tmp_14_9,tmp_14_10,tmp_14_11,tmp_14_12,tmp_14_13,tmp_14_14,1'b0,tmp_14_16,tmp_14_17,tmp_14_18,tmp_14_19,tmp_14_20,tmp_14_21,tmp_14_22,tmp_14_23,tmp_14_24,tmp_14_25,tmp_14_26,tmp_14_27,tmp_14_28,tmp_14_29,tmp_14_30,tmp_14_31};
wire tmp_15_0;
assign tmp_15_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]);
wire tmp_15_1;
assign tmp_15_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]);
wire tmp_15_2;
assign tmp_15_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]);
wire tmp_15_3;
assign tmp_15_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]);
wire tmp_15_4;
assign tmp_15_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]);
wire tmp_15_5;
assign tmp_15_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]);
wire tmp_15_6;
assign tmp_15_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]);
wire tmp_15_7;
assign tmp_15_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]);
wire tmp_15_8;
assign tmp_15_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]);
wire tmp_15_9;
assign tmp_15_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]);
wire tmp_15_10;
assign tmp_15_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]);
wire tmp_15_12;
assign tmp_15_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]);
wire tmp_15_13;
assign tmp_15_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]);
wire tmp_15_14;
assign tmp_15_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]);
wire tmp_15_15;
assign tmp_15_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]);
wire tmp_15_16;
assign tmp_15_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]);
wire tmp_15_17;
assign tmp_15_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]);
wire tmp_15_18;
assign tmp_15_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]);
wire tmp_15_19;
assign tmp_15_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]);
wire tmp_15_20;
assign tmp_15_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]);
wire tmp_15_21;
assign tmp_15_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]);
wire tmp_15_22;
assign tmp_15_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]);
wire tmp_15_23;
assign tmp_15_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]);
wire tmp_15_25;
assign tmp_15_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]);
wire tmp_15_26;
assign tmp_15_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]);
wire tmp_15_27;
assign tmp_15_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]);
wire tmp_15_28;
assign tmp_15_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]);
wire tmp_15_29;
assign tmp_15_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]);
wire tmp_15_30;
assign tmp_15_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]);
wire tmp_15_31;
assign tmp_15_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]);
assign ap_return_15 = {tmp_15_0,tmp_15_1,tmp_15_2,tmp_15_3,tmp_15_4,tmp_15_5,tmp_15_6,tmp_15_7,tmp_15_8,tmp_15_9,tmp_15_10,1'b0,tmp_15_12,tmp_15_13,tmp_15_14,tmp_15_15,tmp_15_16,tmp_15_17,tmp_15_18,tmp_15_19,tmp_15_20,tmp_15_21,tmp_15_22,tmp_15_23,1'b0,tmp_15_25,tmp_15_26,tmp_15_27,tmp_15_28,tmp_15_29,tmp_15_30,tmp_15_31};
wire tmp_16_0;
assign tmp_16_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]);
wire tmp_16_1;
assign tmp_16_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_16_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_16_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_16_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_16_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_16_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_16_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_16_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_16_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_16_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_16_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_16_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_16_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_16_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_16_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_16_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_16_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_16_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_16_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_16_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_16_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_16_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_16_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_16_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_16_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_16_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_16_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_16_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_16_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_16_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_16_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_16_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_16_V_read[1]);
wire tmp_16_2;
assign tmp_16_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_16_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_16_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_16_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_16_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_16_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_16_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_16_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_16_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_16_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_16_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_16_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_16_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_16_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_16_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_16_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_16_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_16_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_16_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_16_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_16_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_16_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_16_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_16_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_16_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_16_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_16_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_16_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_16_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_16_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_16_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_16_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_16_V_read[2]);
wire tmp_16_3;
assign tmp_16_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]);
wire tmp_16_4;
assign tmp_16_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_16_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_16_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_16_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_16_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_16_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_16_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_16_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_16_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_16_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_16_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_16_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_16_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_16_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_16_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_16_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_16_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_16_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_16_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_16_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_16_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_16_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_16_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_16_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_16_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_16_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_16_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_16_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_16_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_16_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_16_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_16_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_16_V_read[4]);
wire tmp_16_6;
assign tmp_16_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_16_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_16_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_16_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_16_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_16_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_16_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_16_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_16_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_16_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_16_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_16_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_16_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_16_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_16_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_16_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_16_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_16_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_16_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_16_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_16_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_16_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_16_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_16_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_16_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_16_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_16_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_16_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_16_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_16_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_16_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_16_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_16_V_read[6]);
wire tmp_16_7;
assign tmp_16_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_16_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_16_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_16_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_16_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_16_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_16_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_16_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_16_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_16_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_16_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_16_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_16_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_16_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_16_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_16_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_16_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_16_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_16_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_16_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_16_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_16_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_16_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_16_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_16_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_16_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_16_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_16_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_16_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_16_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_16_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_16_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_16_V_read[7]);
wire tmp_16_8;
assign tmp_16_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_16_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_16_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_16_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_16_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_16_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_16_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_16_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_16_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_16_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_16_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_16_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_16_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_16_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_16_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_16_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_16_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_16_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_16_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_16_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_16_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_16_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_16_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_16_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_16_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_16_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_16_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_16_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_16_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_16_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_16_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_16_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_16_V_read[8]);
wire tmp_16_9;
assign tmp_16_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_16_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_16_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_16_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_16_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_16_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_16_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_16_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_16_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_16_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_16_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_16_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_16_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_16_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_16_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_16_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_16_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_16_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_16_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_16_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_16_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_16_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_16_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_16_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_16_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_16_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_16_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_16_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_16_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_16_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_16_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_16_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_16_V_read[9]);
wire tmp_16_10;
assign tmp_16_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_16_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_16_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_16_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_16_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_16_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_16_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_16_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_16_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_16_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_16_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_16_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_16_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_16_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_16_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_16_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_16_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_16_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_16_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_16_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_16_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_16_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_16_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_16_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_16_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_16_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_16_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_16_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_16_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_16_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_16_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_16_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_16_V_read[10]);
wire tmp_16_11;
assign tmp_16_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]);
wire tmp_16_13;
assign tmp_16_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_16_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_16_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_16_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_16_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_16_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_16_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_16_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_16_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_16_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_16_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_16_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_16_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_16_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_16_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_16_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_16_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_16_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_16_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_16_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_16_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_16_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_16_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_16_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_16_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_16_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_16_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_16_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_16_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_16_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_16_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_16_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_16_V_read[13]);
wire tmp_16_14;
assign tmp_16_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_16_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_16_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_16_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_16_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_16_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_16_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_16_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_16_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_16_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_16_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_16_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_16_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_16_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_16_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_16_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_16_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_16_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_16_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_16_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_16_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_16_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_16_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_16_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_16_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_16_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_16_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_16_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_16_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_16_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_16_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_16_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_16_V_read[14]);
wire tmp_16_15;
assign tmp_16_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_16_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_16_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_16_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_16_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_16_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_16_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_16_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_16_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_16_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_16_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_16_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_16_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_16_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_16_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_16_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_16_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_16_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_16_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_16_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_16_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_16_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_16_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_16_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_16_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_16_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_16_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_16_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_16_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_16_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_16_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_16_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_16_V_read[15]);
wire tmp_16_16;
assign tmp_16_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_16_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_16_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_16_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_16_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_16_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_16_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_16_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_16_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_16_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_16_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_16_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_16_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_16_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_16_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_16_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_16_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_16_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_16_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_16_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_16_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_16_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_16_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_16_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_16_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_16_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_16_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_16_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_16_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_16_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_16_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_16_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_16_V_read[16]);
wire tmp_16_18;
assign tmp_16_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]);
wire tmp_16_19;
assign tmp_16_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]);
wire tmp_16_20;
assign tmp_16_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_16_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_16_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_16_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_16_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_16_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_16_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_16_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_16_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_16_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_16_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_16_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_16_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_16_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_16_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_16_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_16_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_16_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_16_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_16_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_16_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_16_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_16_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_16_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_16_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_16_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_16_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_16_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_16_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_16_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_16_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_16_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_16_V_read[20]);
wire tmp_16_21;
assign tmp_16_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]);
wire tmp_16_23;
assign tmp_16_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]);
wire tmp_16_24;
assign tmp_16_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]);
wire tmp_16_25;
assign tmp_16_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_16_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_16_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_16_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_16_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_16_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_16_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_16_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_16_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_16_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_16_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_16_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_16_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_16_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_16_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_16_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_16_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_16_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_16_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_16_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_16_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_16_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_16_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_16_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_16_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_16_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_16_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_16_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_16_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_16_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_16_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_16_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_16_V_read[25]);
wire tmp_16_27;
assign tmp_16_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_16_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_16_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_16_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_16_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_16_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_16_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_16_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_16_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_16_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_16_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_16_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_16_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_16_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_16_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_16_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_16_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_16_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_16_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_16_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_16_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_16_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_16_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_16_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_16_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_16_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_16_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_16_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_16_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_16_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_16_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_16_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_16_V_read[27]);
wire tmp_16_28;
assign tmp_16_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_16_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_16_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_16_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_16_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_16_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_16_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_16_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_16_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_16_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_16_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_16_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_16_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_16_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_16_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_16_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_16_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_16_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_16_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_16_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_16_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_16_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_16_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_16_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_16_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_16_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_16_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_16_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_16_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_16_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_16_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_16_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_16_V_read[28]);
wire tmp_16_29;
assign tmp_16_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]);
wire tmp_16_30;
assign tmp_16_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_16_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_16_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_16_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_16_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_16_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_16_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_16_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_16_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_16_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_16_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_16_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_16_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_16_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_16_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_16_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_16_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_16_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_16_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_16_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_16_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_16_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_16_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_16_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_16_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_16_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_16_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_16_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_16_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_16_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_16_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_16_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_16_V_read[30]);
wire tmp_16_31;
assign tmp_16_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]);
assign ap_return_16 = {tmp_16_0,tmp_16_1,tmp_16_2,tmp_16_3,tmp_16_4,1'b0,tmp_16_6,tmp_16_7,tmp_16_8,tmp_16_9,tmp_16_10,tmp_16_11,1'b0,tmp_16_13,tmp_16_14,tmp_16_15,tmp_16_16,1'b0,tmp_16_18,tmp_16_19,tmp_16_20,tmp_16_21,1'b0,tmp_16_23,tmp_16_24,tmp_16_25,1'b0,tmp_16_27,tmp_16_28,tmp_16_29,tmp_16_30,tmp_16_31};
wire tmp_17_0;
assign tmp_17_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]);
wire tmp_17_1;
assign tmp_17_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_17_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_17_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_17_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_17_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_17_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_17_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_17_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_17_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_17_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_17_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_17_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_17_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_17_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_17_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_17_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_17_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_17_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_17_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_17_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_17_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_17_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_17_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_17_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_17_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_17_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_17_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_17_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_17_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_17_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_17_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_17_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_17_V_read[1]);
wire tmp_17_2;
assign tmp_17_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_17_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_17_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_17_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_17_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_17_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_17_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_17_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_17_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_17_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_17_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_17_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_17_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_17_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_17_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_17_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_17_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_17_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_17_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_17_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_17_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_17_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_17_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_17_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_17_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_17_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_17_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_17_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_17_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_17_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_17_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_17_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_17_V_read[2]);
wire tmp_17_3;
assign tmp_17_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]);
wire tmp_17_4;
assign tmp_17_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_17_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_17_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_17_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_17_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_17_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_17_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_17_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_17_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_17_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_17_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_17_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_17_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_17_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_17_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_17_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_17_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_17_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_17_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_17_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_17_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_17_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_17_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_17_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_17_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_17_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_17_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_17_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_17_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_17_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_17_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_17_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_17_V_read[4]);
wire tmp_17_5;
assign tmp_17_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]);
wire tmp_17_6;
assign tmp_17_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_17_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_17_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_17_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_17_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_17_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_17_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_17_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_17_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_17_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_17_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_17_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_17_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_17_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_17_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_17_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_17_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_17_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_17_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_17_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_17_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_17_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_17_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_17_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_17_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_17_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_17_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_17_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_17_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_17_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_17_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_17_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_17_V_read[6]);
wire tmp_17_7;
assign tmp_17_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_17_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_17_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_17_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_17_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_17_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_17_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_17_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_17_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_17_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_17_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_17_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_17_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_17_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_17_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_17_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_17_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_17_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_17_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_17_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_17_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_17_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_17_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_17_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_17_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_17_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_17_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_17_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_17_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_17_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_17_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_17_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_17_V_read[7]);
wire tmp_17_8;
assign tmp_17_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]);
wire tmp_17_9;
assign tmp_17_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_17_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_17_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_17_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_17_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_17_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_17_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_17_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_17_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_17_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_17_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_17_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_17_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_17_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_17_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_17_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_17_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_17_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_17_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_17_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_17_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_17_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_17_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_17_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_17_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_17_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_17_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_17_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_17_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_17_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_17_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_17_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_17_V_read[9]);
wire tmp_17_10;
assign tmp_17_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_17_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_17_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_17_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_17_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_17_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_17_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_17_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_17_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_17_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_17_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_17_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_17_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_17_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_17_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_17_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_17_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_17_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_17_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_17_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_17_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_17_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_17_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_17_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_17_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_17_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_17_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_17_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_17_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_17_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_17_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_17_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_17_V_read[10]);
wire tmp_17_11;
assign tmp_17_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_17_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_17_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_17_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_17_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_17_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_17_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_17_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_17_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_17_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_17_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_17_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_17_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_17_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_17_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_17_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_17_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_17_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_17_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_17_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_17_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_17_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_17_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_17_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_17_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_17_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_17_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_17_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_17_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_17_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_17_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_17_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_17_V_read[11]);
wire tmp_17_12;
assign tmp_17_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_17_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_17_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_17_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_17_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_17_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_17_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_17_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_17_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_17_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_17_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_17_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_17_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_17_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_17_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_17_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_17_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_17_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_17_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_17_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_17_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_17_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_17_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_17_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_17_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_17_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_17_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_17_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_17_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_17_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_17_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_17_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_17_V_read[12]);
wire tmp_17_13;
assign tmp_17_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_17_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_17_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_17_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_17_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_17_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_17_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_17_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_17_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_17_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_17_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_17_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_17_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_17_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_17_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_17_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_17_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_17_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_17_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_17_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_17_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_17_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_17_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_17_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_17_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_17_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_17_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_17_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_17_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_17_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_17_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_17_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_17_V_read[13]);
wire tmp_17_14;
assign tmp_17_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_17_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_17_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_17_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_17_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_17_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_17_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_17_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_17_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_17_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_17_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_17_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_17_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_17_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_17_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_17_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_17_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_17_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_17_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_17_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_17_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_17_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_17_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_17_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_17_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_17_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_17_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_17_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_17_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_17_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_17_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_17_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_17_V_read[14]);
wire tmp_17_15;
assign tmp_17_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_17_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_17_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_17_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_17_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_17_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_17_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_17_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_17_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_17_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_17_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_17_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_17_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_17_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_17_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_17_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_17_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_17_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_17_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_17_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_17_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_17_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_17_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_17_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_17_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_17_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_17_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_17_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_17_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_17_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_17_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_17_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_17_V_read[15]);
wire tmp_17_16;
assign tmp_17_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_17_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_17_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_17_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_17_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_17_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_17_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_17_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_17_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_17_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_17_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_17_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_17_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_17_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_17_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_17_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_17_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_17_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_17_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_17_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_17_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_17_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_17_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_17_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_17_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_17_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_17_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_17_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_17_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_17_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_17_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_17_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_17_V_read[16]);
wire tmp_17_17;
assign tmp_17_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]);
wire tmp_17_18;
assign tmp_17_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_17_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_17_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_17_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_17_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_17_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_17_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_17_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_17_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_17_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_17_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_17_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_17_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_17_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_17_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_17_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_17_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_17_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_17_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_17_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_17_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_17_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_17_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_17_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_17_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_17_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_17_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_17_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_17_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_17_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_17_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_17_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_17_V_read[18]);
wire tmp_17_19;
assign tmp_17_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]);
wire tmp_17_20;
assign tmp_17_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_17_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_17_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_17_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_17_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_17_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_17_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_17_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_17_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_17_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_17_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_17_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_17_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_17_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_17_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_17_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_17_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_17_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_17_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_17_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_17_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_17_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_17_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_17_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_17_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_17_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_17_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_17_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_17_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_17_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_17_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_17_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_17_V_read[20]);
wire tmp_17_21;
assign tmp_17_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]);
wire tmp_17_22;
assign tmp_17_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]);
wire tmp_17_23;
assign tmp_17_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_17_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_17_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_17_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_17_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_17_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_17_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_17_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_17_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_17_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_17_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_17_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_17_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_17_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_17_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_17_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_17_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_17_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_17_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_17_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_17_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_17_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_17_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_17_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_17_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_17_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_17_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_17_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_17_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_17_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_17_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_17_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_17_V_read[23]);
wire tmp_17_24;
assign tmp_17_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_17_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_17_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_17_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_17_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_17_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_17_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_17_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_17_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_17_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_17_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_17_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_17_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_17_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_17_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_17_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_17_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_17_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_17_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_17_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_17_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_17_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_17_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_17_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_17_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_17_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_17_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_17_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_17_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_17_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_17_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_17_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_17_V_read[24]);
wire tmp_17_25;
assign tmp_17_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_17_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_17_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_17_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_17_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_17_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_17_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_17_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_17_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_17_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_17_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_17_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_17_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_17_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_17_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_17_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_17_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_17_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_17_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_17_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_17_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_17_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_17_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_17_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_17_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_17_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_17_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_17_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_17_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_17_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_17_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_17_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_17_V_read[25]);
wire tmp_17_28;
assign tmp_17_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_17_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_17_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_17_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_17_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_17_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_17_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_17_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_17_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_17_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_17_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_17_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_17_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_17_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_17_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_17_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_17_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_17_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_17_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_17_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_17_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_17_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_17_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_17_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_17_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_17_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_17_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_17_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_17_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_17_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_17_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_17_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_17_V_read[28]);
wire tmp_17_29;
assign tmp_17_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_17_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_17_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_17_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_17_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_17_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_17_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_17_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_17_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_17_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_17_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_17_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_17_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_17_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_17_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_17_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_17_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_17_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_17_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_17_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_17_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_17_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_17_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_17_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_17_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_17_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_17_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_17_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_17_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_17_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_17_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_17_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_17_V_read[29]);
wire tmp_17_30;
assign tmp_17_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_17_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_17_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_17_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_17_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_17_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_17_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_17_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_17_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_17_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_17_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_17_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_17_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_17_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_17_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_17_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_17_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_17_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_17_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_17_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_17_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_17_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_17_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_17_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_17_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_17_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_17_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_17_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_17_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_17_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_17_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_17_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_17_V_read[30]);
wire tmp_17_31;
assign tmp_17_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_17_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_17_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_17_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_17_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_17_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_17_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_17_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_17_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_17_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_17_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_17_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_17_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_17_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_17_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_17_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_17_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_17_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_17_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_17_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_17_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_17_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_17_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_17_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_17_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_17_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_17_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_17_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_17_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_17_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_17_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_17_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_17_V_read[31]);
assign ap_return_17 = {tmp_17_0,tmp_17_1,tmp_17_2,tmp_17_3,tmp_17_4,tmp_17_5,tmp_17_6,tmp_17_7,tmp_17_8,tmp_17_9,tmp_17_10,tmp_17_11,tmp_17_12,tmp_17_13,tmp_17_14,tmp_17_15,tmp_17_16,tmp_17_17,tmp_17_18,tmp_17_19,tmp_17_20,tmp_17_21,tmp_17_22,tmp_17_23,tmp_17_24,tmp_17_25,1'b0,1'b0,tmp_17_28,tmp_17_29,tmp_17_30,tmp_17_31};
wire tmp_18_0;
assign tmp_18_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]);
wire tmp_18_1;
assign tmp_18_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_18_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_18_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_18_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_18_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_18_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_18_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_18_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_18_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_18_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_18_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_18_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_18_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_18_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_18_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_18_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_18_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_18_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_18_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_18_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_18_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_18_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_18_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_18_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_18_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_18_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_18_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_18_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_18_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_18_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_18_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_18_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_18_V_read[1]);
wire tmp_18_2;
assign tmp_18_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_18_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_18_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_18_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_18_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_18_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_18_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_18_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_18_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_18_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_18_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_18_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_18_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_18_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_18_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_18_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_18_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_18_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_18_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_18_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_18_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_18_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_18_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_18_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_18_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_18_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_18_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_18_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_18_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_18_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_18_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_18_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_18_V_read[2]);
wire tmp_18_3;
assign tmp_18_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_18_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_18_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_18_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_18_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_18_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_18_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_18_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_18_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_18_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_18_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_18_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_18_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_18_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_18_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_18_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_18_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_18_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_18_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_18_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_18_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_18_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_18_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_18_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_18_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_18_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_18_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_18_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_18_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_18_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_18_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_18_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_18_V_read[3]);
wire tmp_18_4;
assign tmp_18_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_18_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_18_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_18_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_18_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_18_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_18_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_18_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_18_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_18_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_18_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_18_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_18_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_18_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_18_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_18_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_18_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_18_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_18_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_18_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_18_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_18_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_18_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_18_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_18_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_18_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_18_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_18_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_18_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_18_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_18_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_18_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_18_V_read[4]);
wire tmp_18_5;
assign tmp_18_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_18_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_18_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_18_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_18_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_18_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_18_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_18_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_18_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_18_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_18_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_18_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_18_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_18_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_18_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_18_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_18_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_18_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_18_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_18_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_18_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_18_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_18_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_18_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_18_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_18_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_18_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_18_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_18_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_18_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_18_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_18_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_18_V_read[5]);
wire tmp_18_6;
assign tmp_18_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_18_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_18_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_18_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_18_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_18_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_18_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_18_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_18_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_18_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_18_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_18_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_18_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_18_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_18_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_18_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_18_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_18_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_18_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_18_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_18_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_18_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_18_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_18_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_18_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_18_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_18_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_18_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_18_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_18_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_18_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_18_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_18_V_read[6]);
wire tmp_18_7;
assign tmp_18_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]);
wire tmp_18_8;
assign tmp_18_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_18_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_18_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_18_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_18_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_18_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_18_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_18_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_18_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_18_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_18_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_18_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_18_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_18_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_18_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_18_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_18_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_18_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_18_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_18_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_18_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_18_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_18_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_18_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_18_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_18_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_18_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_18_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_18_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_18_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_18_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_18_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_18_V_read[8]);
wire tmp_18_9;
assign tmp_18_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_18_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_18_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_18_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_18_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_18_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_18_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_18_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_18_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_18_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_18_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_18_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_18_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_18_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_18_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_18_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_18_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_18_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_18_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_18_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_18_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_18_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_18_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_18_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_18_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_18_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_18_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_18_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_18_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_18_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_18_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_18_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_18_V_read[9]);
wire tmp_18_10;
assign tmp_18_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]);
wire tmp_18_11;
assign tmp_18_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_18_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_18_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_18_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_18_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_18_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_18_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_18_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_18_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_18_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_18_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_18_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_18_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_18_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_18_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_18_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_18_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_18_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_18_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_18_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_18_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_18_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_18_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_18_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_18_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_18_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_18_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_18_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_18_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_18_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_18_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_18_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_18_V_read[11]);
wire tmp_18_12;
assign tmp_18_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_18_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_18_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_18_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_18_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_18_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_18_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_18_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_18_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_18_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_18_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_18_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_18_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_18_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_18_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_18_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_18_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_18_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_18_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_18_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_18_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_18_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_18_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_18_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_18_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_18_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_18_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_18_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_18_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_18_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_18_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_18_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_18_V_read[12]);
wire tmp_18_13;
assign tmp_18_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_18_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_18_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_18_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_18_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_18_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_18_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_18_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_18_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_18_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_18_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_18_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_18_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_18_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_18_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_18_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_18_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_18_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_18_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_18_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_18_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_18_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_18_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_18_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_18_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_18_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_18_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_18_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_18_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_18_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_18_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_18_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_18_V_read[13]);
wire tmp_18_14;
assign tmp_18_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_18_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_18_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_18_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_18_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_18_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_18_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_18_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_18_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_18_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_18_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_18_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_18_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_18_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_18_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_18_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_18_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_18_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_18_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_18_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_18_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_18_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_18_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_18_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_18_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_18_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_18_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_18_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_18_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_18_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_18_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_18_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_18_V_read[14]);
wire tmp_18_15;
assign tmp_18_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_18_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_18_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_18_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_18_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_18_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_18_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_18_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_18_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_18_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_18_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_18_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_18_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_18_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_18_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_18_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_18_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_18_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_18_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_18_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_18_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_18_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_18_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_18_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_18_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_18_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_18_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_18_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_18_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_18_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_18_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_18_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_18_V_read[15]);
wire tmp_18_16;
assign tmp_18_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]);
wire tmp_18_17;
assign tmp_18_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]);
wire tmp_18_18;
assign tmp_18_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_18_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_18_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_18_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_18_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_18_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_18_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_18_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_18_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_18_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_18_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_18_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_18_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_18_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_18_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_18_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_18_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_18_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_18_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_18_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_18_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_18_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_18_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_18_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_18_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_18_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_18_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_18_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_18_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_18_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_18_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_18_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_18_V_read[18]);
wire tmp_18_19;
assign tmp_18_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]);
wire tmp_18_20;
assign tmp_18_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_18_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_18_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_18_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_18_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_18_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_18_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_18_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_18_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_18_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_18_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_18_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_18_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_18_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_18_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_18_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_18_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_18_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_18_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_18_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_18_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_18_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_18_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_18_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_18_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_18_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_18_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_18_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_18_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_18_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_18_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_18_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_18_V_read[20]);
wire tmp_18_21;
assign tmp_18_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_18_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_18_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_18_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_18_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_18_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_18_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_18_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_18_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_18_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_18_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_18_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_18_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_18_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_18_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_18_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_18_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_18_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_18_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_18_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_18_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_18_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_18_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_18_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_18_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_18_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_18_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_18_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_18_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_18_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_18_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_18_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_18_V_read[21]);
wire tmp_18_22;
assign tmp_18_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_18_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_18_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_18_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_18_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_18_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_18_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_18_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_18_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_18_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_18_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_18_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_18_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_18_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_18_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_18_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_18_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_18_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_18_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_18_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_18_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_18_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_18_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_18_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_18_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_18_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_18_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_18_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_18_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_18_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_18_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_18_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_18_V_read[22]);
wire tmp_18_23;
assign tmp_18_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]);
wire tmp_18_24;
assign tmp_18_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_18_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_18_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_18_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_18_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_18_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_18_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_18_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_18_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_18_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_18_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_18_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_18_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_18_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_18_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_18_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_18_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_18_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_18_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_18_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_18_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_18_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_18_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_18_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_18_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_18_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_18_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_18_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_18_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_18_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_18_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_18_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_18_V_read[24]);
wire tmp_18_25;
assign tmp_18_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]);
wire tmp_18_26;
assign tmp_18_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_18_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_18_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_18_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_18_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_18_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_18_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_18_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_18_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_18_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_18_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_18_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_18_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_18_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_18_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_18_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_18_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_18_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_18_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_18_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_18_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_18_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_18_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_18_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_18_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_18_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_18_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_18_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_18_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_18_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_18_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_18_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_18_V_read[26]);
wire tmp_18_27;
assign tmp_18_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_18_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_18_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_18_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_18_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_18_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_18_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_18_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_18_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_18_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_18_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_18_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_18_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_18_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_18_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_18_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_18_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_18_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_18_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_18_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_18_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_18_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_18_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_18_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_18_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_18_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_18_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_18_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_18_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_18_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_18_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_18_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_18_V_read[27]);
wire tmp_18_28;
assign tmp_18_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_18_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_18_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_18_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_18_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_18_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_18_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_18_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_18_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_18_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_18_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_18_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_18_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_18_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_18_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_18_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_18_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_18_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_18_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_18_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_18_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_18_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_18_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_18_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_18_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_18_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_18_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_18_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_18_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_18_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_18_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_18_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_18_V_read[28]);
wire tmp_18_29;
assign tmp_18_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]);
wire tmp_18_30;
assign tmp_18_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_18_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_18_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_18_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_18_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_18_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_18_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_18_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_18_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_18_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_18_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_18_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_18_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_18_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_18_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_18_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_18_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_18_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_18_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_18_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_18_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_18_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_18_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_18_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_18_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_18_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_18_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_18_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_18_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_18_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_18_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_18_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_18_V_read[30]);
wire tmp_18_31;
assign tmp_18_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]);
assign ap_return_18 = {tmp_18_0,tmp_18_1,tmp_18_2,tmp_18_3,tmp_18_4,tmp_18_5,tmp_18_6,tmp_18_7,tmp_18_8,tmp_18_9,tmp_18_10,tmp_18_11,tmp_18_12,tmp_18_13,tmp_18_14,tmp_18_15,tmp_18_16,tmp_18_17,tmp_18_18,tmp_18_19,tmp_18_20,tmp_18_21,tmp_18_22,tmp_18_23,tmp_18_24,tmp_18_25,tmp_18_26,tmp_18_27,tmp_18_28,tmp_18_29,tmp_18_30,tmp_18_31};
wire tmp_19_0;
assign tmp_19_0 = (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_19_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_19_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_19_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_19_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_19_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_19_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_19_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_19_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_19_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_19_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_19_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_19_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_19_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_19_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_19_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_19_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_19_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_19_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_19_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_19_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_19_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_19_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_19_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_19_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_19_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_19_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_19_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_19_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_19_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_19_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_19_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_19_V_read[0]);
wire tmp_19_1;
assign tmp_19_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_19_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_19_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_19_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_19_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_19_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_19_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_19_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_19_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_19_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_19_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_19_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_19_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_19_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_19_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_19_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_19_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_19_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_19_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_19_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_19_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_19_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_19_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_19_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_19_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_19_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_19_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_19_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_19_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_19_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_19_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_19_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_19_V_read[1]);
wire tmp_19_2;
assign tmp_19_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_19_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_19_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_19_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_19_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_19_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_19_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_19_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_19_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_19_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_19_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_19_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_19_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_19_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_19_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_19_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_19_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_19_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_19_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_19_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_19_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_19_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_19_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_19_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_19_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_19_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_19_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_19_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_19_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_19_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_19_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_19_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_19_V_read[2]);
wire tmp_19_3;
assign tmp_19_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_19_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_19_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_19_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_19_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_19_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_19_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_19_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_19_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_19_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_19_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_19_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_19_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_19_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_19_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_19_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_19_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_19_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_19_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_19_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_19_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_19_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_19_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_19_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_19_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_19_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_19_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_19_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_19_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_19_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_19_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_19_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_19_V_read[3]);
wire tmp_19_4;
assign tmp_19_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_19_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_19_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_19_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_19_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_19_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_19_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_19_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_19_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_19_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_19_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_19_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_19_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_19_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_19_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_19_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_19_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_19_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_19_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_19_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_19_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_19_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_19_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_19_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_19_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_19_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_19_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_19_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_19_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_19_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_19_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_19_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_19_V_read[4]);
wire tmp_19_5;
assign tmp_19_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_19_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_19_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_19_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_19_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_19_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_19_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_19_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_19_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_19_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_19_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_19_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_19_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_19_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_19_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_19_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_19_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_19_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_19_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_19_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_19_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_19_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_19_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_19_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_19_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_19_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_19_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_19_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_19_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_19_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_19_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_19_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_19_V_read[5]);
wire tmp_19_6;
assign tmp_19_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_19_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_19_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_19_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_19_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_19_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_19_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_19_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_19_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_19_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_19_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_19_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_19_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_19_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_19_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_19_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_19_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_19_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_19_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_19_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_19_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_19_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_19_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_19_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_19_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_19_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_19_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_19_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_19_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_19_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_19_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_19_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_19_V_read[6]);
wire tmp_19_7;
assign tmp_19_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]);
wire tmp_19_9;
assign tmp_19_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_19_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_19_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_19_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_19_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_19_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_19_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_19_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_19_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_19_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_19_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_19_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_19_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_19_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_19_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_19_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_19_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_19_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_19_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_19_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_19_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_19_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_19_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_19_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_19_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_19_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_19_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_19_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_19_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_19_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_19_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_19_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_19_V_read[9]);
wire tmp_19_10;
assign tmp_19_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_19_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_19_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_19_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_19_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_19_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_19_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_19_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_19_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_19_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_19_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_19_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_19_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_19_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_19_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_19_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_19_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_19_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_19_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_19_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_19_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_19_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_19_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_19_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_19_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_19_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_19_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_19_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_19_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_19_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_19_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_19_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_19_V_read[10]);
wire tmp_19_11;
assign tmp_19_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_19_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_19_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_19_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_19_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_19_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_19_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_19_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_19_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_19_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_19_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_19_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_19_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_19_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_19_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_19_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_19_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_19_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_19_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_19_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_19_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_19_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_19_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_19_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_19_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_19_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_19_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_19_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_19_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_19_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_19_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_19_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_19_V_read[11]);
wire tmp_19_12;
assign tmp_19_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]);
wire tmp_19_13;
assign tmp_19_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_19_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_19_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_19_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_19_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_19_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_19_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_19_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_19_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_19_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_19_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_19_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_19_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_19_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_19_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_19_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_19_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_19_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_19_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_19_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_19_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_19_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_19_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_19_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_19_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_19_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_19_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_19_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_19_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_19_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_19_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_19_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_19_V_read[13]);
wire tmp_19_14;
assign tmp_19_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_19_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_19_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_19_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_19_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_19_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_19_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_19_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_19_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_19_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_19_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_19_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_19_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_19_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_19_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_19_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_19_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_19_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_19_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_19_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_19_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_19_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_19_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_19_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_19_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_19_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_19_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_19_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_19_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_19_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_19_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_19_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_19_V_read[14]);
wire tmp_19_15;
assign tmp_19_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_19_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_19_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_19_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_19_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_19_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_19_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_19_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_19_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_19_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_19_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_19_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_19_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_19_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_19_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_19_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_19_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_19_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_19_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_19_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_19_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_19_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_19_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_19_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_19_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_19_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_19_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_19_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_19_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_19_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_19_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_19_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_19_V_read[15]);
wire tmp_19_16;
assign tmp_19_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]);
wire tmp_19_17;
assign tmp_19_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_19_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_19_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_19_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_19_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_19_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_19_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_19_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_19_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_19_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_19_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_19_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_19_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_19_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_19_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_19_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_19_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_19_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_19_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_19_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_19_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_19_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_19_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_19_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_19_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_19_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_19_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_19_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_19_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_19_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_19_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_19_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_19_V_read[17]);
wire tmp_19_18;
assign tmp_19_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_19_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_19_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_19_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_19_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_19_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_19_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_19_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_19_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_19_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_19_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_19_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_19_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_19_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_19_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_19_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_19_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_19_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_19_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_19_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_19_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_19_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_19_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_19_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_19_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_19_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_19_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_19_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_19_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_19_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_19_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_19_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_19_V_read[18]);
wire tmp_19_19;
assign tmp_19_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_19_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_19_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_19_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_19_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_19_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_19_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_19_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_19_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_19_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_19_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_19_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_19_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_19_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_19_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_19_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_19_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_19_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_19_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_19_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_19_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_19_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_19_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_19_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_19_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_19_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_19_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_19_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_19_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_19_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_19_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_19_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_19_V_read[19]);
wire tmp_19_20;
assign tmp_19_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_19_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_19_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_19_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_19_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_19_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_19_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_19_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_19_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_19_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_19_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_19_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_19_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_19_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_19_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_19_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_19_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_19_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_19_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_19_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_19_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_19_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_19_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_19_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_19_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_19_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_19_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_19_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_19_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_19_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_19_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_19_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_19_V_read[20]);
wire tmp_19_21;
assign tmp_19_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_19_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_19_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_19_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_19_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_19_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_19_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_19_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_19_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_19_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_19_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_19_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_19_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_19_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_19_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_19_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_19_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_19_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_19_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_19_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_19_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_19_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_19_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_19_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_19_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_19_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_19_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_19_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_19_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_19_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_19_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_19_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_19_V_read[21]);
wire tmp_19_22;
assign tmp_19_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]);
wire tmp_19_23;
assign tmp_19_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_19_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_19_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_19_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_19_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_19_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_19_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_19_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_19_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_19_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_19_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_19_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_19_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_19_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_19_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_19_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_19_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_19_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_19_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_19_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_19_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_19_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_19_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_19_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_19_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_19_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_19_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_19_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_19_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_19_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_19_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_19_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_19_V_read[23]);
wire tmp_19_24;
assign tmp_19_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_19_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_19_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_19_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_19_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_19_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_19_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_19_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_19_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_19_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_19_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_19_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_19_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_19_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_19_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_19_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_19_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_19_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_19_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_19_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_19_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_19_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_19_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_19_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_19_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_19_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_19_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_19_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_19_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_19_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_19_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_19_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_19_V_read[24]);
wire tmp_19_25;
assign tmp_19_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_19_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_19_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_19_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_19_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_19_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_19_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_19_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_19_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_19_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_19_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_19_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_19_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_19_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_19_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_19_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_19_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_19_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_19_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_19_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_19_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_19_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_19_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_19_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_19_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_19_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_19_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_19_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_19_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_19_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_19_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_19_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_19_V_read[25]);
wire tmp_19_27;
assign tmp_19_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_19_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_19_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_19_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_19_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_19_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_19_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_19_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_19_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_19_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_19_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_19_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_19_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_19_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_19_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_19_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_19_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_19_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_19_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_19_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_19_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_19_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_19_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_19_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_19_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_19_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_19_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_19_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_19_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_19_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_19_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_19_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_19_V_read[27]);
wire tmp_19_28;
assign tmp_19_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_19_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_19_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_19_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_19_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_19_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_19_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_19_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_19_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_19_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_19_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_19_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_19_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_19_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_19_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_19_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_19_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_19_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_19_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_19_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_19_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_19_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_19_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_19_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_19_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_19_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_19_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_19_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_19_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_19_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_19_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_19_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_19_V_read[28]);
wire tmp_19_29;
assign tmp_19_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_19_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_19_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_19_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_19_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_19_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_19_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_19_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_19_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_19_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_19_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_19_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_19_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_19_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_19_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_19_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_19_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_19_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_19_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_19_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_19_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_19_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_19_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_19_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_19_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_19_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_19_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_19_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_19_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_19_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_19_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_19_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_19_V_read[29]);
assign ap_return_19 = {tmp_19_0,tmp_19_1,tmp_19_2,tmp_19_3,tmp_19_4,tmp_19_5,tmp_19_6,tmp_19_7,1'b0,tmp_19_9,tmp_19_10,tmp_19_11,tmp_19_12,tmp_19_13,tmp_19_14,tmp_19_15,tmp_19_16,tmp_19_17,tmp_19_18,tmp_19_19,tmp_19_20,tmp_19_21,tmp_19_22,tmp_19_23,tmp_19_24,tmp_19_25,1'b0,tmp_19_27,tmp_19_28,tmp_19_29,1'b0,1'b0};
wire tmp_20_0;
assign tmp_20_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]);
wire tmp_20_1;
assign tmp_20_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_20_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_20_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_20_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_20_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_20_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_20_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_20_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_20_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_20_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_20_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_20_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_20_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_20_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_20_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_20_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_20_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_20_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_20_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_20_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_20_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_20_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_20_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_20_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_20_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_20_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_20_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_20_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_20_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_20_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_20_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_20_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_20_V_read[1]);
wire tmp_20_3;
assign tmp_20_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]);
wire tmp_20_4;
assign tmp_20_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_20_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_20_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_20_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_20_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_20_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_20_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_20_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_20_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_20_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_20_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_20_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_20_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_20_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_20_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_20_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_20_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_20_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_20_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_20_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_20_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_20_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_20_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_20_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_20_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_20_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_20_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_20_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_20_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_20_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_20_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_20_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_20_V_read[4]);
wire tmp_20_5;
assign tmp_20_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]);
wire tmp_20_6;
assign tmp_20_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_20_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_20_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_20_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_20_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_20_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_20_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_20_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_20_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_20_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_20_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_20_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_20_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_20_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_20_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_20_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_20_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_20_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_20_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_20_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_20_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_20_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_20_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_20_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_20_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_20_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_20_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_20_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_20_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_20_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_20_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_20_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_20_V_read[6]);
wire tmp_20_7;
assign tmp_20_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_20_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_20_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_20_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_20_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_20_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_20_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_20_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_20_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_20_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_20_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_20_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_20_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_20_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_20_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_20_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_20_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_20_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_20_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_20_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_20_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_20_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_20_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_20_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_20_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_20_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_20_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_20_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_20_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_20_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_20_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_20_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_20_V_read[7]);
wire tmp_20_8;
assign tmp_20_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]);
wire tmp_20_9;
assign tmp_20_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_20_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_20_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_20_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_20_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_20_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_20_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_20_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_20_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_20_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_20_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_20_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_20_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_20_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_20_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_20_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_20_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_20_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_20_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_20_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_20_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_20_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_20_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_20_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_20_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_20_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_20_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_20_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_20_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_20_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_20_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_20_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_20_V_read[9]);
wire tmp_20_10;
assign tmp_20_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_20_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_20_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_20_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_20_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_20_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_20_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_20_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_20_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_20_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_20_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_20_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_20_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_20_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_20_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_20_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_20_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_20_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_20_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_20_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_20_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_20_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_20_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_20_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_20_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_20_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_20_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_20_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_20_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_20_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_20_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_20_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_20_V_read[10]);
wire tmp_20_11;
assign tmp_20_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_20_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_20_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_20_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_20_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_20_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_20_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_20_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_20_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_20_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_20_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_20_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_20_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_20_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_20_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_20_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_20_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_20_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_20_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_20_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_20_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_20_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_20_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_20_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_20_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_20_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_20_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_20_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_20_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_20_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_20_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_20_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_20_V_read[11]);
wire tmp_20_13;
assign tmp_20_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_20_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_20_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_20_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_20_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_20_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_20_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_20_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_20_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_20_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_20_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_20_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_20_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_20_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_20_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_20_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_20_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_20_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_20_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_20_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_20_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_20_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_20_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_20_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_20_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_20_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_20_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_20_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_20_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_20_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_20_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_20_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_20_V_read[13]);
wire tmp_20_14;
assign tmp_20_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_20_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_20_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_20_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_20_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_20_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_20_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_20_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_20_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_20_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_20_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_20_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_20_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_20_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_20_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_20_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_20_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_20_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_20_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_20_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_20_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_20_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_20_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_20_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_20_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_20_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_20_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_20_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_20_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_20_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_20_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_20_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_20_V_read[14]);
wire tmp_20_16;
assign tmp_20_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]);
wire tmp_20_17;
assign tmp_20_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]);
wire tmp_20_18;
assign tmp_20_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_20_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_20_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_20_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_20_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_20_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_20_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_20_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_20_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_20_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_20_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_20_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_20_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_20_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_20_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_20_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_20_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_20_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_20_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_20_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_20_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_20_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_20_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_20_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_20_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_20_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_20_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_20_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_20_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_20_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_20_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_20_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_20_V_read[18]);
wire tmp_20_20;
assign tmp_20_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_20_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_20_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_20_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_20_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_20_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_20_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_20_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_20_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_20_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_20_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_20_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_20_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_20_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_20_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_20_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_20_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_20_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_20_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_20_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_20_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_20_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_20_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_20_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_20_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_20_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_20_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_20_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_20_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_20_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_20_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_20_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_20_V_read[20]);
wire tmp_20_21;
assign tmp_20_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]);
wire tmp_20_22;
assign tmp_20_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_20_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_20_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_20_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_20_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_20_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_20_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_20_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_20_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_20_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_20_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_20_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_20_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_20_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_20_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_20_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_20_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_20_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_20_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_20_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_20_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_20_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_20_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_20_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_20_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_20_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_20_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_20_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_20_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_20_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_20_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_20_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_20_V_read[22]);
wire tmp_20_23;
assign tmp_20_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_20_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_20_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_20_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_20_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_20_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_20_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_20_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_20_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_20_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_20_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_20_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_20_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_20_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_20_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_20_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_20_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_20_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_20_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_20_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_20_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_20_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_20_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_20_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_20_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_20_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_20_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_20_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_20_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_20_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_20_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_20_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_20_V_read[23]);
wire tmp_20_24;
assign tmp_20_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_20_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_20_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_20_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_20_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_20_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_20_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_20_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_20_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_20_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_20_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_20_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_20_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_20_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_20_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_20_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_20_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_20_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_20_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_20_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_20_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_20_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_20_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_20_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_20_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_20_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_20_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_20_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_20_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_20_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_20_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_20_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_20_V_read[24]);
wire tmp_20_25;
assign tmp_20_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_20_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_20_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_20_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_20_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_20_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_20_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_20_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_20_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_20_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_20_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_20_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_20_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_20_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_20_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_20_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_20_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_20_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_20_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_20_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_20_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_20_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_20_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_20_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_20_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_20_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_20_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_20_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_20_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_20_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_20_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_20_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_20_V_read[25]);
wire tmp_20_26;
assign tmp_20_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_20_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_20_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_20_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_20_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_20_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_20_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_20_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_20_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_20_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_20_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_20_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_20_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_20_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_20_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_20_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_20_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_20_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_20_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_20_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_20_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_20_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_20_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_20_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_20_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_20_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_20_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_20_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_20_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_20_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_20_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_20_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_20_V_read[26]);
wire tmp_20_27;
assign tmp_20_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_20_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_20_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_20_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_20_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_20_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_20_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_20_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_20_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_20_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_20_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_20_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_20_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_20_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_20_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_20_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_20_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_20_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_20_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_20_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_20_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_20_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_20_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_20_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_20_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_20_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_20_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_20_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_20_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_20_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_20_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_20_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_20_V_read[27]);
wire tmp_20_28;
assign tmp_20_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]);
wire tmp_20_29;
assign tmp_20_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_20_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_20_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_20_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_20_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_20_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_20_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_20_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_20_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_20_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_20_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_20_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_20_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_20_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_20_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_20_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_20_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_20_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_20_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_20_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_20_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_20_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_20_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_20_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_20_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_20_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_20_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_20_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_20_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_20_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_20_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_20_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_20_V_read[29]);
wire tmp_20_30;
assign tmp_20_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_20_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_20_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_20_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_20_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_20_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_20_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_20_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_20_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_20_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_20_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_20_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_20_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_20_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_20_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_20_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_20_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_20_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_20_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_20_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_20_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_20_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_20_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_20_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_20_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_20_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_20_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_20_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_20_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_20_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_20_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_20_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_20_V_read[30]);
wire tmp_20_31;
assign tmp_20_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_20_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_20_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_20_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_20_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_20_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_20_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_20_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_20_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_20_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_20_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_20_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_20_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_20_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_20_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_20_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_20_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_20_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_20_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_20_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_20_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_20_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_20_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_20_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_20_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_20_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_20_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_20_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_20_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_20_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_20_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_20_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_20_V_read[31]);
assign ap_return_20 = {tmp_20_0,tmp_20_1,1'b0,tmp_20_3,tmp_20_4,tmp_20_5,tmp_20_6,tmp_20_7,tmp_20_8,tmp_20_9,tmp_20_10,tmp_20_11,1'b0,tmp_20_13,tmp_20_14,1'b0,tmp_20_16,tmp_20_17,tmp_20_18,1'b0,tmp_20_20,tmp_20_21,tmp_20_22,tmp_20_23,tmp_20_24,tmp_20_25,tmp_20_26,tmp_20_27,tmp_20_28,tmp_20_29,tmp_20_30,tmp_20_31};
wire tmp_21_0;
assign tmp_21_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]);
wire tmp_21_1;
assign tmp_21_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_21_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_21_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_21_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_21_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_21_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_21_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_21_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_21_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_21_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_21_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_21_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_21_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_21_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_21_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_21_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_21_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_21_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_21_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_21_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_21_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_21_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_21_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_21_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_21_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_21_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_21_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_21_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_21_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_21_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_21_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_21_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_21_V_read[1]);
wire tmp_21_2;
assign tmp_21_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_21_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_21_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_21_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_21_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_21_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_21_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_21_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_21_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_21_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_21_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_21_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_21_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_21_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_21_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_21_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_21_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_21_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_21_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_21_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_21_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_21_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_21_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_21_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_21_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_21_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_21_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_21_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_21_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_21_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_21_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_21_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_21_V_read[2]);
wire tmp_21_3;
assign tmp_21_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_21_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_21_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_21_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_21_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_21_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_21_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_21_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_21_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_21_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_21_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_21_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_21_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_21_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_21_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_21_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_21_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_21_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_21_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_21_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_21_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_21_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_21_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_21_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_21_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_21_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_21_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_21_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_21_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_21_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_21_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_21_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_21_V_read[3]);
wire tmp_21_4;
assign tmp_21_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_21_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_21_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_21_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_21_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_21_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_21_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_21_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_21_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_21_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_21_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_21_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_21_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_21_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_21_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_21_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_21_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_21_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_21_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_21_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_21_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_21_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_21_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_21_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_21_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_21_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_21_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_21_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_21_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_21_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_21_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_21_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_21_V_read[4]);
wire tmp_21_5;
assign tmp_21_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_21_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_21_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_21_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_21_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_21_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_21_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_21_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_21_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_21_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_21_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_21_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_21_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_21_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_21_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_21_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_21_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_21_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_21_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_21_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_21_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_21_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_21_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_21_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_21_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_21_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_21_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_21_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_21_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_21_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_21_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_21_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_21_V_read[5]);
wire tmp_21_6;
assign tmp_21_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_21_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_21_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_21_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_21_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_21_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_21_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_21_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_21_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_21_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_21_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_21_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_21_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_21_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_21_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_21_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_21_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_21_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_21_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_21_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_21_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_21_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_21_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_21_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_21_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_21_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_21_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_21_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_21_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_21_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_21_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_21_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_21_V_read[6]);
wire tmp_21_7;
assign tmp_21_7 = (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]);
wire tmp_21_9;
assign tmp_21_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_21_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_21_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_21_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_21_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_21_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_21_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_21_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_21_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_21_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_21_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_21_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_21_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_21_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_21_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_21_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_21_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_21_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_21_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_21_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_21_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_21_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_21_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_21_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_21_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_21_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_21_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_21_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_21_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_21_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_21_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_21_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_21_V_read[9]);
wire tmp_21_10;
assign tmp_21_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_21_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_21_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_21_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_21_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_21_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_21_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_21_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_21_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_21_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_21_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_21_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_21_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_21_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_21_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_21_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_21_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_21_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_21_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_21_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_21_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_21_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_21_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_21_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_21_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_21_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_21_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_21_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_21_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_21_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_21_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_21_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_21_V_read[10]);
wire tmp_21_11;
assign tmp_21_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_21_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_21_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_21_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_21_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_21_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_21_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_21_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_21_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_21_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_21_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_21_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_21_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_21_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_21_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_21_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_21_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_21_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_21_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_21_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_21_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_21_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_21_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_21_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_21_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_21_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_21_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_21_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_21_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_21_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_21_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_21_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_21_V_read[11]);
wire tmp_21_12;
assign tmp_21_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_21_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_21_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_21_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_21_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_21_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_21_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_21_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_21_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_21_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_21_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_21_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_21_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_21_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_21_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_21_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_21_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_21_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_21_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_21_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_21_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_21_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_21_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_21_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_21_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_21_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_21_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_21_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_21_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_21_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_21_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_21_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_21_V_read[12]);
wire tmp_21_13;
assign tmp_21_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_21_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_21_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_21_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_21_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_21_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_21_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_21_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_21_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_21_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_21_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_21_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_21_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_21_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_21_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_21_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_21_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_21_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_21_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_21_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_21_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_21_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_21_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_21_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_21_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_21_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_21_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_21_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_21_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_21_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_21_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_21_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_21_V_read[13]);
wire tmp_21_14;
assign tmp_21_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_21_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_21_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_21_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_21_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_21_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_21_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_21_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_21_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_21_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_21_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_21_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_21_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_21_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_21_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_21_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_21_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_21_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_21_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_21_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_21_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_21_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_21_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_21_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_21_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_21_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_21_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_21_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_21_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_21_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_21_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_21_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_21_V_read[14]);
wire tmp_21_16;
assign tmp_21_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]);
wire tmp_21_17;
assign tmp_21_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_21_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_21_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_21_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_21_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_21_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_21_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_21_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_21_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_21_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_21_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_21_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_21_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_21_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_21_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_21_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_21_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_21_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_21_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_21_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_21_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_21_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_21_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_21_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_21_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_21_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_21_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_21_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_21_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_21_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_21_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_21_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_21_V_read[17]);
wire tmp_21_18;
assign tmp_21_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_21_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_21_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_21_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_21_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_21_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_21_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_21_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_21_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_21_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_21_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_21_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_21_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_21_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_21_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_21_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_21_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_21_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_21_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_21_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_21_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_21_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_21_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_21_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_21_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_21_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_21_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_21_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_21_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_21_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_21_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_21_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_21_V_read[18]);
wire tmp_21_20;
assign tmp_21_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_21_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_21_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_21_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_21_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_21_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_21_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_21_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_21_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_21_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_21_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_21_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_21_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_21_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_21_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_21_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_21_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_21_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_21_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_21_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_21_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_21_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_21_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_21_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_21_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_21_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_21_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_21_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_21_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_21_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_21_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_21_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_21_V_read[20]);
wire tmp_21_21;
assign tmp_21_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]);
wire tmp_21_22;
assign tmp_21_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_21_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_21_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_21_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_21_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_21_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_21_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_21_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_21_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_21_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_21_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_21_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_21_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_21_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_21_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_21_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_21_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_21_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_21_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_21_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_21_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_21_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_21_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_21_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_21_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_21_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_21_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_21_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_21_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_21_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_21_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_21_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_21_V_read[22]);
wire tmp_21_23;
assign tmp_21_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_21_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_21_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_21_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_21_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_21_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_21_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_21_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_21_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_21_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_21_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_21_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_21_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_21_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_21_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_21_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_21_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_21_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_21_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_21_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_21_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_21_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_21_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_21_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_21_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_21_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_21_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_21_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_21_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_21_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_21_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_21_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_21_V_read[23]);
wire tmp_21_24;
assign tmp_21_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]);
wire tmp_21_25;
assign tmp_21_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_21_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_21_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_21_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_21_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_21_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_21_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_21_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_21_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_21_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_21_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_21_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_21_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_21_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_21_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_21_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_21_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_21_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_21_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_21_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_21_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_21_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_21_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_21_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_21_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_21_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_21_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_21_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_21_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_21_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_21_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_21_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_21_V_read[25]);
wire tmp_21_26;
assign tmp_21_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]);
wire tmp_21_27;
assign tmp_21_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_21_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_21_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_21_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_21_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_21_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_21_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_21_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_21_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_21_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_21_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_21_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_21_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_21_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_21_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_21_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_21_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_21_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_21_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_21_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_21_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_21_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_21_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_21_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_21_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_21_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_21_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_21_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_21_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_21_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_21_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_21_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_21_V_read[27]);
wire tmp_21_28;
assign tmp_21_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]);
wire tmp_21_29;
assign tmp_21_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]);
wire tmp_21_30;
assign tmp_21_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]);
wire tmp_21_31;
assign tmp_21_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]);
assign ap_return_21 = {tmp_21_0,tmp_21_1,tmp_21_2,tmp_21_3,tmp_21_4,tmp_21_5,tmp_21_6,tmp_21_7,1'b0,tmp_21_9,tmp_21_10,tmp_21_11,tmp_21_12,tmp_21_13,tmp_21_14,1'b0,tmp_21_16,tmp_21_17,tmp_21_18,1'b0,tmp_21_20,tmp_21_21,tmp_21_22,tmp_21_23,tmp_21_24,tmp_21_25,tmp_21_26,tmp_21_27,tmp_21_28,tmp_21_29,tmp_21_30,tmp_21_31};
wire tmp_22_0;
assign tmp_22_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]);
wire tmp_22_1;
assign tmp_22_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]);
wire tmp_22_2;
assign tmp_22_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_22_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_22_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_22_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_22_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_22_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_22_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_22_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_22_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_22_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_22_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_22_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_22_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_22_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_22_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_22_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_22_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_22_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_22_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_22_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_22_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_22_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_22_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_22_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_22_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_22_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_22_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_22_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_22_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_22_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_22_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_22_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_22_V_read[2]);
wire tmp_22_3;
assign tmp_22_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]);
wire tmp_22_4;
assign tmp_22_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_22_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_22_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_22_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_22_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_22_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_22_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_22_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_22_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_22_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_22_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_22_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_22_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_22_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_22_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_22_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_22_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_22_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_22_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_22_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_22_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_22_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_22_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_22_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_22_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_22_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_22_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_22_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_22_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_22_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_22_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_22_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_22_V_read[4]);
wire tmp_22_6;
assign tmp_22_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]);
wire tmp_22_7;
assign tmp_22_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_22_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_22_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_22_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_22_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_22_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_22_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_22_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_22_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_22_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_22_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_22_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_22_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_22_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_22_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_22_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_22_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_22_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_22_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_22_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_22_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_22_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_22_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_22_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_22_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_22_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_22_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_22_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_22_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_22_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_22_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_22_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_22_V_read[7]);
wire tmp_22_8;
assign tmp_22_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]);
wire tmp_22_9;
assign tmp_22_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_22_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_22_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_22_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_22_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_22_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_22_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_22_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_22_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_22_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_22_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_22_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_22_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_22_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_22_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_22_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_22_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_22_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_22_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_22_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_22_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_22_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_22_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_22_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_22_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_22_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_22_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_22_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_22_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_22_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_22_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_22_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_22_V_read[9]);
wire tmp_22_10;
assign tmp_22_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_22_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_22_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_22_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_22_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_22_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_22_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_22_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_22_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_22_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_22_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_22_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_22_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_22_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_22_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_22_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_22_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_22_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_22_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_22_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_22_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_22_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_22_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_22_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_22_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_22_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_22_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_22_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_22_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_22_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_22_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_22_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_22_V_read[10]);
wire tmp_22_11;
assign tmp_22_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_22_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_22_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_22_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_22_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_22_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_22_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_22_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_22_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_22_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_22_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_22_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_22_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_22_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_22_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_22_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_22_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_22_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_22_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_22_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_22_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_22_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_22_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_22_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_22_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_22_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_22_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_22_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_22_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_22_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_22_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_22_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_22_V_read[11]);
wire tmp_22_12;
assign tmp_22_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_22_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_22_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_22_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_22_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_22_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_22_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_22_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_22_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_22_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_22_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_22_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_22_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_22_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_22_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_22_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_22_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_22_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_22_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_22_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_22_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_22_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_22_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_22_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_22_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_22_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_22_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_22_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_22_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_22_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_22_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_22_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_22_V_read[12]);
wire tmp_22_13;
assign tmp_22_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_22_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_22_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_22_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_22_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_22_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_22_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_22_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_22_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_22_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_22_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_22_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_22_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_22_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_22_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_22_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_22_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_22_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_22_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_22_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_22_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_22_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_22_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_22_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_22_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_22_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_22_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_22_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_22_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_22_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_22_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_22_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_22_V_read[13]);
wire tmp_22_14;
assign tmp_22_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_22_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_22_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_22_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_22_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_22_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_22_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_22_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_22_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_22_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_22_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_22_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_22_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_22_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_22_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_22_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_22_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_22_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_22_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_22_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_22_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_22_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_22_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_22_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_22_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_22_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_22_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_22_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_22_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_22_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_22_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_22_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_22_V_read[14]);
wire tmp_22_15;
assign tmp_22_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_22_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_22_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_22_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_22_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_22_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_22_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_22_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_22_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_22_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_22_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_22_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_22_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_22_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_22_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_22_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_22_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_22_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_22_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_22_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_22_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_22_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_22_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_22_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_22_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_22_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_22_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_22_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_22_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_22_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_22_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_22_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_22_V_read[15]);
wire tmp_22_17;
assign tmp_22_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]);
wire tmp_22_18;
assign tmp_22_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_22_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_22_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_22_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_22_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_22_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_22_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_22_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_22_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_22_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_22_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_22_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_22_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_22_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_22_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_22_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_22_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_22_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_22_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_22_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_22_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_22_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_22_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_22_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_22_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_22_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_22_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_22_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_22_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_22_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_22_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_22_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_22_V_read[18]);
wire tmp_22_20;
assign tmp_22_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_22_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_22_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_22_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_22_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_22_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_22_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_22_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_22_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_22_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_22_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_22_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_22_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_22_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_22_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_22_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_22_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_22_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_22_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_22_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_22_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_22_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_22_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_22_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_22_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_22_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_22_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_22_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_22_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_22_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_22_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_22_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_22_V_read[20]);
wire tmp_22_21;
assign tmp_22_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]);
wire tmp_22_22;
assign tmp_22_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]);
wire tmp_22_23;
assign tmp_22_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]);
wire tmp_22_24;
assign tmp_22_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_22_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_22_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_22_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_22_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_22_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_22_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_22_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_22_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_22_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_22_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_22_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_22_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_22_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_22_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_22_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_22_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_22_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_22_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_22_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_22_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_22_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_22_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_22_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_22_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_22_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_22_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_22_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_22_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_22_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_22_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_22_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_22_V_read[24]);
wire tmp_22_25;
assign tmp_22_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_22_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_22_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_22_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_22_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_22_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_22_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_22_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_22_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_22_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_22_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_22_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_22_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_22_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_22_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_22_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_22_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_22_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_22_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_22_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_22_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_22_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_22_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_22_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_22_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_22_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_22_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_22_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_22_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_22_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_22_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_22_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_22_V_read[25]);
wire tmp_22_26;
assign tmp_22_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]);
wire tmp_22_27;
assign tmp_22_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_22_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_22_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_22_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_22_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_22_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_22_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_22_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_22_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_22_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_22_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_22_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_22_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_22_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_22_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_22_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_22_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_22_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_22_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_22_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_22_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_22_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_22_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_22_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_22_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_22_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_22_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_22_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_22_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_22_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_22_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_22_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_22_V_read[27]);
wire tmp_22_28;
assign tmp_22_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_22_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_22_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_22_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_22_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_22_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_22_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_22_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_22_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_22_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_22_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_22_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_22_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_22_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_22_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_22_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_22_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_22_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_22_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_22_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_22_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_22_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_22_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_22_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_22_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_22_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_22_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_22_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_22_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_22_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_22_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_22_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_22_V_read[28]);
wire tmp_22_29;
assign tmp_22_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]);
wire tmp_22_30;
assign tmp_22_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_22_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_22_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_22_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_22_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_22_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_22_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_22_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_22_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_22_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_22_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_22_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_22_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_22_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_22_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_22_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_22_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_22_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_22_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_22_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_22_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_22_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_22_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_22_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_22_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_22_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_22_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_22_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_22_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_22_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_22_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_22_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_22_V_read[30]);
wire tmp_22_31;
assign tmp_22_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]);
assign ap_return_22 = {tmp_22_0,tmp_22_1,tmp_22_2,tmp_22_3,tmp_22_4,1'b0,tmp_22_6,tmp_22_7,tmp_22_8,tmp_22_9,tmp_22_10,tmp_22_11,tmp_22_12,tmp_22_13,tmp_22_14,tmp_22_15,1'b0,tmp_22_17,tmp_22_18,1'b0,tmp_22_20,tmp_22_21,tmp_22_22,tmp_22_23,tmp_22_24,tmp_22_25,tmp_22_26,tmp_22_27,tmp_22_28,tmp_22_29,tmp_22_30,tmp_22_31};
wire tmp_23_0;
assign tmp_23_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]);
wire tmp_23_1;
assign tmp_23_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]);
wire tmp_23_2;
assign tmp_23_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_23_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_23_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_23_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_23_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_23_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_23_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_23_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_23_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_23_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_23_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_23_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_23_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_23_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_23_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_23_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_23_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_23_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_23_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_23_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_23_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_23_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_23_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_23_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_23_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_23_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_23_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_23_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_23_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_23_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_23_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_23_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_23_V_read[2]);
wire tmp_23_3;
assign tmp_23_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_23_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_23_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_23_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_23_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_23_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_23_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_23_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_23_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_23_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_23_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_23_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_23_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_23_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_23_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_23_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_23_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_23_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_23_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_23_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_23_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_23_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_23_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_23_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_23_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_23_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_23_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_23_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_23_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_23_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_23_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_23_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_23_V_read[3]);
wire tmp_23_4;
assign tmp_23_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_23_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_23_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_23_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_23_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_23_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_23_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_23_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_23_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_23_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_23_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_23_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_23_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_23_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_23_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_23_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_23_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_23_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_23_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_23_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_23_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_23_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_23_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_23_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_23_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_23_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_23_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_23_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_23_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_23_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_23_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_23_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_23_V_read[4]);
wire tmp_23_5;
assign tmp_23_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_23_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_23_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_23_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_23_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_23_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_23_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_23_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_23_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_23_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_23_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_23_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_23_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_23_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_23_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_23_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_23_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_23_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_23_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_23_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_23_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_23_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_23_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_23_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_23_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_23_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_23_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_23_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_23_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_23_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_23_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_23_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_23_V_read[5]);
wire tmp_23_6;
assign tmp_23_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_23_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_23_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_23_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_23_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_23_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_23_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_23_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_23_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_23_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_23_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_23_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_23_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_23_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_23_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_23_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_23_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_23_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_23_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_23_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_23_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_23_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_23_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_23_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_23_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_23_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_23_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_23_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_23_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_23_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_23_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_23_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_23_V_read[6]);
wire tmp_23_8;
assign tmp_23_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_23_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_23_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_23_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_23_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_23_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_23_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_23_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_23_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_23_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_23_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_23_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_23_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_23_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_23_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_23_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_23_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_23_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_23_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_23_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_23_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_23_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_23_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_23_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_23_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_23_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_23_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_23_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_23_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_23_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_23_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_23_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_23_V_read[8]);
wire tmp_23_9;
assign tmp_23_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_23_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_23_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_23_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_23_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_23_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_23_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_23_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_23_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_23_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_23_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_23_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_23_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_23_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_23_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_23_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_23_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_23_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_23_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_23_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_23_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_23_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_23_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_23_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_23_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_23_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_23_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_23_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_23_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_23_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_23_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_23_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_23_V_read[9]);
wire tmp_23_10;
assign tmp_23_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_23_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_23_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_23_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_23_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_23_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_23_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_23_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_23_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_23_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_23_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_23_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_23_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_23_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_23_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_23_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_23_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_23_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_23_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_23_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_23_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_23_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_23_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_23_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_23_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_23_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_23_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_23_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_23_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_23_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_23_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_23_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_23_V_read[10]);
wire tmp_23_11;
assign tmp_23_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_23_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_23_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_23_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_23_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_23_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_23_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_23_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_23_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_23_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_23_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_23_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_23_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_23_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_23_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_23_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_23_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_23_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_23_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_23_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_23_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_23_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_23_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_23_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_23_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_23_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_23_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_23_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_23_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_23_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_23_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_23_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_23_V_read[11]);
wire tmp_23_12;
assign tmp_23_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_23_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_23_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_23_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_23_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_23_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_23_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_23_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_23_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_23_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_23_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_23_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_23_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_23_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_23_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_23_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_23_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_23_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_23_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_23_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_23_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_23_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_23_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_23_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_23_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_23_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_23_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_23_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_23_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_23_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_23_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_23_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_23_V_read[12]);
wire tmp_23_13;
assign tmp_23_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_23_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_23_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_23_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_23_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_23_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_23_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_23_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_23_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_23_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_23_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_23_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_23_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_23_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_23_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_23_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_23_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_23_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_23_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_23_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_23_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_23_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_23_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_23_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_23_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_23_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_23_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_23_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_23_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_23_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_23_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_23_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_23_V_read[13]);
wire tmp_23_14;
assign tmp_23_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_23_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_23_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_23_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_23_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_23_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_23_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_23_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_23_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_23_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_23_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_23_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_23_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_23_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_23_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_23_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_23_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_23_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_23_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_23_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_23_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_23_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_23_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_23_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_23_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_23_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_23_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_23_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_23_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_23_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_23_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_23_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_23_V_read[14]);
wire tmp_23_15;
assign tmp_23_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]);
wire tmp_23_16;
assign tmp_23_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_23_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_23_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_23_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_23_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_23_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_23_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_23_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_23_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_23_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_23_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_23_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_23_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_23_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_23_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_23_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_23_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_23_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_23_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_23_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_23_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_23_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_23_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_23_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_23_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_23_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_23_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_23_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_23_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_23_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_23_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_23_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_23_V_read[16]);
wire tmp_23_17;
assign tmp_23_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]);
wire tmp_23_18;
assign tmp_23_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]);
wire tmp_23_19;
assign tmp_23_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_23_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_23_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_23_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_23_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_23_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_23_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_23_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_23_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_23_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_23_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_23_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_23_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_23_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_23_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_23_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_23_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_23_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_23_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_23_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_23_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_23_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_23_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_23_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_23_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_23_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_23_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_23_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_23_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_23_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_23_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_23_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_23_V_read[19]);
wire tmp_23_20;
assign tmp_23_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_23_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_23_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_23_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_23_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_23_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_23_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_23_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_23_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_23_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_23_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_23_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_23_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_23_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_23_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_23_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_23_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_23_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_23_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_23_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_23_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_23_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_23_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_23_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_23_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_23_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_23_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_23_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_23_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_23_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_23_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_23_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_23_V_read[20]);
wire tmp_23_21;
assign tmp_23_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_23_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_23_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_23_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_23_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_23_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_23_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_23_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_23_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_23_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_23_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_23_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_23_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_23_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_23_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_23_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_23_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_23_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_23_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_23_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_23_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_23_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_23_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_23_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_23_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_23_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_23_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_23_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_23_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_23_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_23_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_23_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_23_V_read[21]);
wire tmp_23_22;
assign tmp_23_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_23_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_23_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_23_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_23_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_23_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_23_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_23_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_23_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_23_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_23_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_23_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_23_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_23_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_23_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_23_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_23_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_23_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_23_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_23_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_23_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_23_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_23_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_23_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_23_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_23_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_23_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_23_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_23_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_23_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_23_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_23_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_23_V_read[22]);
wire tmp_23_23;
assign tmp_23_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_23_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_23_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_23_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_23_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_23_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_23_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_23_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_23_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_23_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_23_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_23_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_23_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_23_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_23_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_23_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_23_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_23_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_23_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_23_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_23_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_23_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_23_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_23_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_23_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_23_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_23_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_23_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_23_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_23_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_23_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_23_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_23_V_read[23]);
wire tmp_23_24;
assign tmp_23_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_23_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_23_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_23_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_23_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_23_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_23_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_23_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_23_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_23_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_23_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_23_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_23_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_23_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_23_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_23_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_23_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_23_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_23_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_23_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_23_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_23_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_23_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_23_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_23_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_23_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_23_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_23_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_23_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_23_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_23_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_23_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_23_V_read[24]);
wire tmp_23_26;
assign tmp_23_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]);
wire tmp_23_27;
assign tmp_23_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_23_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_23_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_23_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_23_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_23_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_23_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_23_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_23_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_23_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_23_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_23_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_23_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_23_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_23_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_23_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_23_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_23_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_23_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_23_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_23_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_23_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_23_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_23_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_23_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_23_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_23_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_23_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_23_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_23_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_23_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_23_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_23_V_read[27]);
wire tmp_23_28;
assign tmp_23_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_23_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_23_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_23_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_23_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_23_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_23_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_23_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_23_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_23_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_23_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_23_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_23_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_23_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_23_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_23_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_23_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_23_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_23_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_23_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_23_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_23_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_23_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_23_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_23_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_23_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_23_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_23_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_23_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_23_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_23_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_23_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_23_V_read[28]);
wire tmp_23_29;
assign tmp_23_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]);
wire tmp_23_30;
assign tmp_23_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_23_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_23_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_23_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_23_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_23_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_23_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_23_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_23_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_23_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_23_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_23_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_23_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_23_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_23_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_23_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_23_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_23_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_23_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_23_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_23_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_23_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_23_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_23_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_23_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_23_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_23_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_23_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_23_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_23_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_23_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_23_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_23_V_read[30]);
wire tmp_23_31;
assign tmp_23_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_23_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_23_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_23_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_23_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_23_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_23_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_23_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_23_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_23_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_23_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_23_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_23_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_23_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_23_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_23_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_23_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_23_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_23_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_23_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_23_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_23_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_23_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_23_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_23_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_23_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_23_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_23_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_23_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_23_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_23_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_23_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_23_V_read[31]);
assign ap_return_23 = {tmp_23_0,tmp_23_1,tmp_23_2,tmp_23_3,tmp_23_4,tmp_23_5,tmp_23_6,1'b0,tmp_23_8,tmp_23_9,tmp_23_10,tmp_23_11,tmp_23_12,tmp_23_13,tmp_23_14,tmp_23_15,tmp_23_16,tmp_23_17,tmp_23_18,tmp_23_19,tmp_23_20,tmp_23_21,tmp_23_22,tmp_23_23,tmp_23_24,1'b0,tmp_23_26,tmp_23_27,tmp_23_28,tmp_23_29,tmp_23_30,tmp_23_31};
wire tmp_24_0;
assign tmp_24_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]);
wire tmp_24_1;
assign tmp_24_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_24_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_24_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_24_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_24_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_24_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_24_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_24_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_24_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_24_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_24_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_24_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_24_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_24_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_24_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_24_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_24_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_24_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_24_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_24_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_24_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_24_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_24_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_24_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_24_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_24_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_24_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_24_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_24_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_24_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_24_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_24_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_24_V_read[1]);
wire tmp_24_2;
assign tmp_24_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_24_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_24_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_24_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_24_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_24_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_24_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_24_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_24_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_24_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_24_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_24_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_24_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_24_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_24_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_24_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_24_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_24_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_24_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_24_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_24_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_24_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_24_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_24_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_24_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_24_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_24_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_24_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_24_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_24_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_24_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_24_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_24_V_read[2]);
wire tmp_24_3;
assign tmp_24_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_24_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_24_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_24_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_24_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_24_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_24_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_24_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_24_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_24_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_24_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_24_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_24_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_24_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_24_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_24_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_24_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_24_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_24_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_24_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_24_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_24_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_24_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_24_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_24_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_24_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_24_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_24_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_24_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_24_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_24_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_24_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_24_V_read[3]);
wire tmp_24_4;
assign tmp_24_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_24_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_24_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_24_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_24_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_24_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_24_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_24_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_24_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_24_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_24_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_24_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_24_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_24_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_24_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_24_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_24_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_24_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_24_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_24_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_24_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_24_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_24_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_24_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_24_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_24_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_24_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_24_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_24_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_24_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_24_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_24_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_24_V_read[4]);
wire tmp_24_6;
assign tmp_24_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_24_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_24_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_24_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_24_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_24_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_24_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_24_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_24_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_24_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_24_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_24_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_24_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_24_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_24_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_24_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_24_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_24_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_24_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_24_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_24_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_24_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_24_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_24_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_24_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_24_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_24_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_24_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_24_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_24_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_24_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_24_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_24_V_read[6]);
wire tmp_24_7;
assign tmp_24_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_24_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_24_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_24_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_24_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_24_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_24_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_24_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_24_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_24_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_24_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_24_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_24_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_24_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_24_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_24_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_24_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_24_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_24_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_24_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_24_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_24_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_24_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_24_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_24_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_24_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_24_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_24_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_24_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_24_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_24_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_24_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_24_V_read[7]);
wire tmp_24_8;
assign tmp_24_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]);
wire tmp_24_9;
assign tmp_24_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_24_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_24_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_24_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_24_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_24_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_24_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_24_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_24_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_24_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_24_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_24_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_24_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_24_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_24_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_24_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_24_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_24_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_24_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_24_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_24_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_24_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_24_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_24_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_24_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_24_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_24_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_24_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_24_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_24_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_24_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_24_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_24_V_read[9]);
wire tmp_24_10;
assign tmp_24_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_24_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_24_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_24_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_24_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_24_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_24_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_24_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_24_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_24_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_24_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_24_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_24_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_24_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_24_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_24_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_24_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_24_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_24_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_24_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_24_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_24_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_24_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_24_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_24_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_24_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_24_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_24_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_24_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_24_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_24_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_24_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_24_V_read[10]);
wire tmp_24_11;
assign tmp_24_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_24_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_24_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_24_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_24_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_24_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_24_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_24_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_24_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_24_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_24_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_24_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_24_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_24_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_24_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_24_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_24_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_24_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_24_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_24_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_24_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_24_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_24_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_24_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_24_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_24_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_24_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_24_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_24_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_24_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_24_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_24_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_24_V_read[11]);
wire tmp_24_12;
assign tmp_24_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_24_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_24_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_24_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_24_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_24_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_24_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_24_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_24_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_24_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_24_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_24_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_24_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_24_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_24_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_24_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_24_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_24_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_24_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_24_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_24_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_24_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_24_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_24_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_24_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_24_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_24_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_24_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_24_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_24_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_24_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_24_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_24_V_read[12]);
wire tmp_24_13;
assign tmp_24_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_24_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_24_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_24_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_24_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_24_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_24_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_24_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_24_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_24_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_24_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_24_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_24_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_24_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_24_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_24_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_24_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_24_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_24_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_24_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_24_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_24_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_24_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_24_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_24_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_24_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_24_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_24_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_24_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_24_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_24_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_24_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_24_V_read[13]);
wire tmp_24_14;
assign tmp_24_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_24_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_24_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_24_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_24_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_24_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_24_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_24_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_24_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_24_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_24_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_24_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_24_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_24_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_24_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_24_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_24_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_24_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_24_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_24_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_24_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_24_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_24_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_24_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_24_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_24_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_24_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_24_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_24_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_24_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_24_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_24_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_24_V_read[14]);
wire tmp_24_15;
assign tmp_24_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_24_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_24_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_24_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_24_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_24_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_24_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_24_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_24_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_24_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_24_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_24_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_24_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_24_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_24_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_24_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_24_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_24_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_24_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_24_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_24_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_24_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_24_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_24_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_24_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_24_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_24_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_24_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_24_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_24_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_24_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_24_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_24_V_read[15]);
wire tmp_24_16;
assign tmp_24_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]);
wire tmp_24_17;
assign tmp_24_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_24_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_24_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_24_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_24_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_24_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_24_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_24_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_24_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_24_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_24_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_24_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_24_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_24_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_24_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_24_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_24_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_24_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_24_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_24_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_24_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_24_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_24_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_24_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_24_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_24_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_24_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_24_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_24_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_24_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_24_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_24_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_24_V_read[17]);
wire tmp_24_18;
assign tmp_24_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_24_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_24_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_24_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_24_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_24_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_24_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_24_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_24_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_24_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_24_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_24_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_24_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_24_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_24_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_24_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_24_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_24_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_24_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_24_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_24_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_24_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_24_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_24_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_24_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_24_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_24_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_24_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_24_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_24_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_24_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_24_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_24_V_read[18]);
wire tmp_24_19;
assign tmp_24_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_24_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_24_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_24_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_24_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_24_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_24_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_24_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_24_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_24_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_24_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_24_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_24_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_24_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_24_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_24_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_24_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_24_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_24_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_24_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_24_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_24_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_24_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_24_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_24_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_24_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_24_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_24_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_24_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_24_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_24_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_24_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_24_V_read[19]);
wire tmp_24_20;
assign tmp_24_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_24_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_24_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_24_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_24_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_24_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_24_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_24_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_24_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_24_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_24_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_24_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_24_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_24_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_24_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_24_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_24_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_24_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_24_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_24_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_24_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_24_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_24_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_24_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_24_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_24_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_24_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_24_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_24_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_24_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_24_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_24_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_24_V_read[20]);
wire tmp_24_21;
assign tmp_24_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_24_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_24_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_24_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_24_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_24_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_24_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_24_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_24_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_24_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_24_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_24_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_24_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_24_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_24_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_24_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_24_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_24_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_24_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_24_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_24_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_24_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_24_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_24_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_24_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_24_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_24_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_24_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_24_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_24_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_24_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_24_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_24_V_read[21]);
wire tmp_24_22;
assign tmp_24_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_24_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_24_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_24_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_24_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_24_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_24_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_24_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_24_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_24_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_24_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_24_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_24_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_24_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_24_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_24_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_24_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_24_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_24_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_24_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_24_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_24_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_24_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_24_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_24_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_24_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_24_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_24_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_24_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_24_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_24_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_24_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_24_V_read[22]);
wire tmp_24_23;
assign tmp_24_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]);
wire tmp_24_24;
assign tmp_24_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_24_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_24_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_24_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_24_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_24_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_24_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_24_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_24_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_24_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_24_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_24_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_24_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_24_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_24_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_24_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_24_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_24_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_24_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_24_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_24_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_24_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_24_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_24_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_24_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_24_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_24_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_24_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_24_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_24_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_24_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_24_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_24_V_read[24]);
wire tmp_24_25;
assign tmp_24_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_24_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_24_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_24_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_24_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_24_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_24_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_24_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_24_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_24_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_24_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_24_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_24_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_24_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_24_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_24_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_24_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_24_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_24_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_24_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_24_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_24_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_24_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_24_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_24_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_24_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_24_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_24_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_24_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_24_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_24_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_24_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_24_V_read[25]);
wire tmp_24_27;
assign tmp_24_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]);
wire tmp_24_28;
assign tmp_24_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_24_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_24_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_24_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_24_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_24_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_24_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_24_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_24_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_24_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_24_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_24_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_24_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_24_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_24_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_24_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_24_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_24_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_24_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_24_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_24_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_24_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_24_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_24_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_24_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_24_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_24_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_24_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_24_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_24_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_24_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_24_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_24_V_read[28]);
wire tmp_24_29;
assign tmp_24_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]);
wire tmp_24_30;
assign tmp_24_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_24_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_24_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_24_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_24_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_24_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_24_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_24_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_24_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_24_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_24_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_24_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_24_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_24_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_24_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_24_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_24_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_24_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_24_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_24_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_24_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_24_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_24_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_24_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_24_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_24_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_24_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_24_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_24_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_24_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_24_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_24_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_24_V_read[30]);
wire tmp_24_31;
assign tmp_24_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]);
assign ap_return_24 = {tmp_24_0,tmp_24_1,tmp_24_2,tmp_24_3,tmp_24_4,1'b0,tmp_24_6,tmp_24_7,tmp_24_8,tmp_24_9,tmp_24_10,tmp_24_11,tmp_24_12,tmp_24_13,tmp_24_14,tmp_24_15,tmp_24_16,tmp_24_17,tmp_24_18,tmp_24_19,tmp_24_20,tmp_24_21,tmp_24_22,tmp_24_23,tmp_24_24,tmp_24_25,1'b0,tmp_24_27,tmp_24_28,tmp_24_29,tmp_24_30,tmp_24_31};
wire tmp_25_0;
assign tmp_25_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_25_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_25_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_25_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_25_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_25_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_25_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_25_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_25_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_25_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_25_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_25_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_25_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_25_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_25_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_25_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_25_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_25_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_25_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_25_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_25_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_25_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_25_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_25_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_25_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_25_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_25_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_25_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_25_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_25_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_25_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_25_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_25_V_read[0]);
wire tmp_25_1;
assign tmp_25_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_25_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_25_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_25_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_25_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_25_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_25_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_25_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_25_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_25_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_25_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_25_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_25_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_25_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_25_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_25_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_25_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_25_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_25_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_25_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_25_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_25_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_25_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_25_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_25_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_25_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_25_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_25_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_25_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_25_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_25_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_25_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_25_V_read[1]);
wire tmp_25_2;
assign tmp_25_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_25_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_25_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_25_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_25_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_25_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_25_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_25_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_25_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_25_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_25_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_25_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_25_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_25_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_25_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_25_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_25_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_25_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_25_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_25_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_25_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_25_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_25_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_25_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_25_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_25_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_25_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_25_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_25_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_25_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_25_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_25_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_25_V_read[2]);
wire tmp_25_3;
assign tmp_25_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_25_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_25_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_25_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_25_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_25_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_25_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_25_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_25_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_25_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_25_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_25_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_25_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_25_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_25_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_25_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_25_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_25_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_25_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_25_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_25_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_25_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_25_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_25_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_25_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_25_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_25_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_25_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_25_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_25_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_25_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_25_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_25_V_read[3]);
wire tmp_25_4;
assign tmp_25_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_25_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_25_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_25_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_25_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_25_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_25_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_25_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_25_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_25_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_25_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_25_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_25_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_25_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_25_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_25_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_25_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_25_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_25_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_25_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_25_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_25_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_25_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_25_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_25_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_25_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_25_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_25_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_25_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_25_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_25_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_25_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_25_V_read[4]);
wire tmp_25_6;
assign tmp_25_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_25_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_25_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_25_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_25_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_25_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_25_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_25_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_25_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_25_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_25_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_25_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_25_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_25_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_25_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_25_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_25_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_25_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_25_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_25_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_25_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_25_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_25_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_25_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_25_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_25_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_25_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_25_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_25_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_25_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_25_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_25_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_25_V_read[6]);
wire tmp_25_7;
assign tmp_25_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_25_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_25_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_25_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_25_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_25_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_25_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_25_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_25_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_25_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_25_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_25_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_25_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_25_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_25_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_25_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_25_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_25_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_25_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_25_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_25_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_25_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_25_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_25_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_25_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_25_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_25_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_25_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_25_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_25_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_25_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_25_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_25_V_read[7]);
wire tmp_25_8;
assign tmp_25_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]);
wire tmp_25_9;
assign tmp_25_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_25_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_25_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_25_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_25_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_25_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_25_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_25_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_25_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_25_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_25_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_25_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_25_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_25_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_25_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_25_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_25_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_25_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_25_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_25_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_25_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_25_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_25_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_25_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_25_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_25_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_25_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_25_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_25_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_25_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_25_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_25_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_25_V_read[9]);
wire tmp_25_10;
assign tmp_25_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_25_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_25_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_25_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_25_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_25_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_25_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_25_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_25_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_25_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_25_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_25_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_25_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_25_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_25_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_25_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_25_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_25_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_25_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_25_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_25_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_25_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_25_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_25_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_25_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_25_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_25_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_25_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_25_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_25_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_25_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_25_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_25_V_read[10]);
wire tmp_25_11;
assign tmp_25_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_25_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_25_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_25_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_25_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_25_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_25_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_25_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_25_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_25_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_25_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_25_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_25_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_25_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_25_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_25_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_25_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_25_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_25_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_25_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_25_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_25_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_25_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_25_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_25_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_25_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_25_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_25_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_25_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_25_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_25_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_25_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_25_V_read[11]);
wire tmp_25_12;
assign tmp_25_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_25_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_25_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_25_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_25_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_25_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_25_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_25_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_25_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_25_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_25_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_25_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_25_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_25_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_25_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_25_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_25_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_25_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_25_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_25_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_25_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_25_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_25_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_25_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_25_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_25_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_25_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_25_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_25_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_25_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_25_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_25_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_25_V_read[12]);
wire tmp_25_13;
assign tmp_25_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]);
wire tmp_25_14;
assign tmp_25_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_25_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_25_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_25_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_25_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_25_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_25_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_25_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_25_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_25_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_25_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_25_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_25_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_25_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_25_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_25_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_25_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_25_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_25_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_25_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_25_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_25_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_25_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_25_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_25_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_25_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_25_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_25_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_25_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_25_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_25_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_25_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_25_V_read[14]);
wire tmp_25_15;
assign tmp_25_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_25_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_25_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_25_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_25_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_25_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_25_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_25_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_25_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_25_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_25_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_25_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_25_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_25_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_25_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_25_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_25_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_25_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_25_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_25_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_25_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_25_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_25_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_25_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_25_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_25_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_25_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_25_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_25_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_25_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_25_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_25_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_25_V_read[15]);
wire tmp_25_16;
assign tmp_25_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_25_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_25_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_25_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_25_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_25_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_25_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_25_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_25_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_25_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_25_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_25_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_25_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_25_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_25_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_25_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_25_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_25_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_25_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_25_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_25_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_25_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_25_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_25_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_25_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_25_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_25_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_25_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_25_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_25_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_25_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_25_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_25_V_read[16]);
wire tmp_25_17;
assign tmp_25_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_25_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_25_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_25_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_25_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_25_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_25_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_25_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_25_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_25_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_25_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_25_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_25_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_25_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_25_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_25_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_25_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_25_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_25_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_25_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_25_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_25_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_25_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_25_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_25_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_25_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_25_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_25_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_25_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_25_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_25_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_25_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_25_V_read[17]);
wire tmp_25_18;
assign tmp_25_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_25_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_25_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_25_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_25_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_25_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_25_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_25_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_25_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_25_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_25_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_25_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_25_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_25_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_25_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_25_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_25_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_25_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_25_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_25_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_25_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_25_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_25_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_25_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_25_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_25_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_25_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_25_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_25_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_25_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_25_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_25_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_25_V_read[18]);
wire tmp_25_19;
assign tmp_25_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_25_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_25_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_25_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_25_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_25_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_25_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_25_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_25_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_25_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_25_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_25_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_25_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_25_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_25_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_25_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_25_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_25_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_25_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_25_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_25_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_25_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_25_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_25_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_25_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_25_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_25_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_25_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_25_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_25_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_25_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_25_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_25_V_read[19]);
wire tmp_25_20;
assign tmp_25_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_25_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_25_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_25_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_25_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_25_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_25_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_25_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_25_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_25_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_25_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_25_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_25_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_25_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_25_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_25_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_25_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_25_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_25_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_25_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_25_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_25_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_25_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_25_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_25_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_25_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_25_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_25_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_25_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_25_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_25_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_25_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_25_V_read[20]);
wire tmp_25_21;
assign tmp_25_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]);
wire tmp_25_22;
assign tmp_25_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_25_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_25_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_25_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_25_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_25_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_25_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_25_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_25_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_25_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_25_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_25_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_25_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_25_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_25_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_25_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_25_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_25_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_25_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_25_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_25_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_25_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_25_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_25_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_25_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_25_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_25_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_25_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_25_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_25_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_25_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_25_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_25_V_read[22]);
wire tmp_25_24;
assign tmp_25_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]);
wire tmp_25_25;
assign tmp_25_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_25_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_25_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_25_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_25_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_25_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_25_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_25_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_25_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_25_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_25_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_25_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_25_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_25_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_25_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_25_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_25_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_25_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_25_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_25_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_25_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_25_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_25_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_25_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_25_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_25_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_25_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_25_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_25_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_25_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_25_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_25_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_25_V_read[25]);
wire tmp_25_26;
assign tmp_25_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_25_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_25_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_25_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_25_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_25_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_25_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_25_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_25_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_25_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_25_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_25_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_25_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_25_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_25_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_25_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_25_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_25_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_25_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_25_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_25_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_25_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_25_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_25_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_25_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_25_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_25_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_25_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_25_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_25_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_25_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_25_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_25_V_read[26]);
wire tmp_25_27;
assign tmp_25_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_25_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_25_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_25_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_25_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_25_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_25_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_25_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_25_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_25_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_25_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_25_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_25_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_25_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_25_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_25_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_25_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_25_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_25_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_25_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_25_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_25_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_25_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_25_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_25_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_25_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_25_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_25_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_25_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_25_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_25_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_25_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_25_V_read[27]);
wire tmp_25_28;
assign tmp_25_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_25_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_25_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_25_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_25_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_25_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_25_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_25_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_25_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_25_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_25_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_25_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_25_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_25_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_25_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_25_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_25_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_25_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_25_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_25_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_25_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_25_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_25_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_25_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_25_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_25_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_25_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_25_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_25_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_25_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_25_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_25_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_25_V_read[28]);
wire tmp_25_30;
assign tmp_25_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_25_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_25_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_25_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_25_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_25_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_25_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_25_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_25_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_25_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_25_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_25_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_25_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_25_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_25_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_25_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_25_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_25_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_25_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_25_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_25_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_25_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_25_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_25_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_25_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_25_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_25_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_25_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_25_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_25_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_25_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_25_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_25_V_read[30]);
assign ap_return_25 = {tmp_25_0,tmp_25_1,tmp_25_2,tmp_25_3,tmp_25_4,1'b0,tmp_25_6,tmp_25_7,tmp_25_8,tmp_25_9,tmp_25_10,tmp_25_11,tmp_25_12,tmp_25_13,tmp_25_14,tmp_25_15,tmp_25_16,tmp_25_17,tmp_25_18,tmp_25_19,tmp_25_20,tmp_25_21,tmp_25_22,1'b0,tmp_25_24,tmp_25_25,tmp_25_26,tmp_25_27,tmp_25_28,1'b0,tmp_25_30,1'b0};
wire tmp_26_0;
assign tmp_26_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_26_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_26_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_26_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_26_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_26_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_26_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_26_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_26_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_26_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_26_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_26_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_26_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_26_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_26_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_26_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_26_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_26_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_26_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_26_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_26_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_26_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_26_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_26_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_26_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_26_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_26_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_26_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_26_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_26_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_26_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_26_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_26_V_read[0]);
wire tmp_26_1;
assign tmp_26_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_26_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_26_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_26_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_26_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_26_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_26_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_26_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_26_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_26_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_26_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_26_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_26_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_26_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_26_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_26_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_26_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_26_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_26_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_26_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_26_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_26_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_26_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_26_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_26_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_26_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_26_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_26_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_26_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_26_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_26_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_26_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_26_V_read[1]);
wire tmp_26_2;
assign tmp_26_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]);
wire tmp_26_3;
assign tmp_26_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_26_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_26_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_26_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_26_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_26_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_26_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_26_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_26_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_26_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_26_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_26_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_26_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_26_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_26_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_26_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_26_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_26_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_26_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_26_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_26_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_26_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_26_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_26_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_26_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_26_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_26_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_26_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_26_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_26_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_26_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_26_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_26_V_read[3]);
wire tmp_26_4;
assign tmp_26_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_26_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_26_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_26_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_26_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_26_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_26_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_26_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_26_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_26_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_26_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_26_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_26_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_26_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_26_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_26_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_26_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_26_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_26_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_26_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_26_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_26_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_26_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_26_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_26_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_26_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_26_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_26_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_26_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_26_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_26_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_26_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_26_V_read[4]);
wire tmp_26_5;
assign tmp_26_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_26_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_26_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_26_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_26_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_26_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_26_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_26_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_26_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_26_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_26_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_26_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_26_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_26_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_26_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_26_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_26_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_26_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_26_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_26_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_26_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_26_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_26_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_26_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_26_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_26_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_26_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_26_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_26_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_26_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_26_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_26_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_26_V_read[5]);
wire tmp_26_6;
assign tmp_26_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_26_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_26_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_26_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_26_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_26_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_26_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_26_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_26_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_26_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_26_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_26_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_26_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_26_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_26_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_26_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_26_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_26_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_26_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_26_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_26_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_26_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_26_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_26_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_26_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_26_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_26_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_26_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_26_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_26_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_26_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_26_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_26_V_read[6]);
wire tmp_26_7;
assign tmp_26_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_26_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_26_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_26_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_26_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_26_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_26_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_26_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_26_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_26_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_26_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_26_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_26_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_26_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_26_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_26_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_26_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_26_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_26_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_26_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_26_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_26_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_26_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_26_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_26_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_26_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_26_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_26_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_26_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_26_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_26_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_26_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_26_V_read[7]);
wire tmp_26_8;
assign tmp_26_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_26_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_26_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_26_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_26_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_26_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_26_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_26_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_26_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_26_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_26_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_26_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_26_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_26_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_26_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_26_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_26_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_26_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_26_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_26_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_26_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_26_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_26_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_26_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_26_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_26_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_26_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_26_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_26_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_26_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_26_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_26_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_26_V_read[8]);
wire tmp_26_9;
assign tmp_26_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]);
wire tmp_26_10;
assign tmp_26_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_26_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_26_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_26_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_26_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_26_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_26_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_26_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_26_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_26_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_26_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_26_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_26_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_26_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_26_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_26_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_26_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_26_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_26_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_26_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_26_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_26_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_26_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_26_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_26_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_26_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_26_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_26_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_26_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_26_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_26_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_26_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_26_V_read[10]);
wire tmp_26_11;
assign tmp_26_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_26_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_26_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_26_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_26_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_26_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_26_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_26_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_26_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_26_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_26_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_26_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_26_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_26_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_26_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_26_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_26_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_26_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_26_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_26_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_26_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_26_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_26_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_26_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_26_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_26_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_26_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_26_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_26_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_26_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_26_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_26_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_26_V_read[11]);
wire tmp_26_12;
assign tmp_26_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_26_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_26_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_26_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_26_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_26_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_26_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_26_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_26_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_26_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_26_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_26_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_26_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_26_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_26_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_26_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_26_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_26_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_26_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_26_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_26_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_26_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_26_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_26_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_26_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_26_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_26_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_26_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_26_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_26_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_26_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_26_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_26_V_read[12]);
wire tmp_26_13;
assign tmp_26_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_26_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_26_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_26_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_26_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_26_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_26_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_26_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_26_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_26_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_26_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_26_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_26_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_26_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_26_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_26_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_26_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_26_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_26_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_26_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_26_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_26_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_26_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_26_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_26_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_26_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_26_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_26_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_26_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_26_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_26_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_26_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_26_V_read[13]);
wire tmp_26_14;
assign tmp_26_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_26_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_26_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_26_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_26_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_26_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_26_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_26_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_26_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_26_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_26_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_26_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_26_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_26_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_26_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_26_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_26_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_26_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_26_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_26_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_26_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_26_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_26_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_26_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_26_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_26_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_26_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_26_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_26_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_26_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_26_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_26_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_26_V_read[14]);
wire tmp_26_15;
assign tmp_26_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_26_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_26_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_26_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_26_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_26_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_26_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_26_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_26_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_26_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_26_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_26_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_26_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_26_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_26_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_26_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_26_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_26_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_26_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_26_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_26_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_26_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_26_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_26_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_26_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_26_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_26_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_26_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_26_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_26_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_26_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_26_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_26_V_read[15]);
wire tmp_26_16;
assign tmp_26_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]);
wire tmp_26_17;
assign tmp_26_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]);
wire tmp_26_18;
assign tmp_26_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_26_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_26_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_26_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_26_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_26_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_26_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_26_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_26_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_26_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_26_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_26_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_26_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_26_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_26_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_26_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_26_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_26_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_26_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_26_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_26_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_26_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_26_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_26_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_26_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_26_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_26_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_26_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_26_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_26_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_26_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_26_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_26_V_read[18]);
wire tmp_26_19;
assign tmp_26_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_26_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_26_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_26_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_26_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_26_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_26_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_26_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_26_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_26_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_26_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_26_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_26_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_26_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_26_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_26_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_26_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_26_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_26_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_26_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_26_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_26_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_26_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_26_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_26_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_26_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_26_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_26_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_26_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_26_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_26_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_26_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_26_V_read[19]);
wire tmp_26_20;
assign tmp_26_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_26_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_26_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_26_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_26_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_26_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_26_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_26_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_26_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_26_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_26_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_26_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_26_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_26_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_26_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_26_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_26_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_26_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_26_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_26_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_26_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_26_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_26_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_26_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_26_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_26_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_26_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_26_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_26_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_26_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_26_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_26_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_26_V_read[20]);
wire tmp_26_23;
assign tmp_26_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]);
wire tmp_26_24;
assign tmp_26_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]);
wire tmp_26_25;
assign tmp_26_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_26_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_26_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_26_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_26_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_26_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_26_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_26_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_26_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_26_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_26_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_26_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_26_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_26_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_26_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_26_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_26_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_26_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_26_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_26_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_26_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_26_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_26_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_26_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_26_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_26_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_26_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_26_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_26_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_26_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_26_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_26_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_26_V_read[25]);
wire tmp_26_26;
assign tmp_26_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_26_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_26_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_26_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_26_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_26_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_26_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_26_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_26_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_26_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_26_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_26_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_26_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_26_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_26_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_26_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_26_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_26_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_26_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_26_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_26_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_26_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_26_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_26_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_26_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_26_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_26_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_26_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_26_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_26_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_26_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_26_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_26_V_read[26]);
wire tmp_26_27;
assign tmp_26_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_26_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_26_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_26_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_26_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_26_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_26_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_26_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_26_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_26_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_26_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_26_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_26_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_26_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_26_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_26_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_26_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_26_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_26_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_26_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_26_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_26_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_26_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_26_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_26_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_26_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_26_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_26_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_26_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_26_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_26_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_26_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_26_V_read[27]);
wire tmp_26_28;
assign tmp_26_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_26_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_26_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_26_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_26_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_26_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_26_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_26_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_26_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_26_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_26_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_26_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_26_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_26_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_26_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_26_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_26_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_26_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_26_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_26_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_26_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_26_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_26_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_26_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_26_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_26_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_26_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_26_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_26_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_26_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_26_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_26_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_26_V_read[28]);
wire tmp_26_29;
assign tmp_26_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]);
wire tmp_26_30;
assign tmp_26_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_26_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_26_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_26_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_26_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_26_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_26_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_26_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_26_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_26_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_26_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_26_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_26_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_26_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_26_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_26_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_26_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_26_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_26_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_26_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_26_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_26_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_26_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_26_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_26_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_26_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_26_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_26_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_26_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_26_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_26_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_26_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_26_V_read[30]);
wire tmp_26_31;
assign tmp_26_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_26_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_26_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_26_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_26_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_26_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_26_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_26_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_26_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_26_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_26_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_26_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_26_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_26_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_26_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_26_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_26_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_26_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_26_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_26_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_26_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_26_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_26_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_26_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_26_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_26_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_26_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_26_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_26_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_26_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_26_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_26_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_26_V_read[31]);
assign ap_return_26 = {tmp_26_0,tmp_26_1,tmp_26_2,tmp_26_3,tmp_26_4,tmp_26_5,tmp_26_6,tmp_26_7,tmp_26_8,tmp_26_9,tmp_26_10,tmp_26_11,tmp_26_12,tmp_26_13,tmp_26_14,tmp_26_15,tmp_26_16,tmp_26_17,tmp_26_18,tmp_26_19,tmp_26_20,1'b0,1'b0,tmp_26_23,tmp_26_24,tmp_26_25,tmp_26_26,tmp_26_27,tmp_26_28,tmp_26_29,tmp_26_30,tmp_26_31};
wire tmp_27_0;
assign tmp_27_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_27_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_27_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_27_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_27_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_27_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_27_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_27_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_27_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_27_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_27_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_27_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_27_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_27_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_27_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_27_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_27_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_27_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_27_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_27_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_27_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_27_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_27_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_27_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_27_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_27_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_27_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_27_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_27_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_27_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_27_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_27_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_27_V_read[0]);
wire tmp_27_1;
assign tmp_27_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_27_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_27_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_27_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_27_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_27_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_27_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_27_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_27_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_27_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_27_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_27_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_27_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_27_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_27_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_27_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_27_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_27_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_27_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_27_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_27_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_27_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_27_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_27_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_27_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_27_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_27_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_27_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_27_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_27_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_27_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_27_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_27_V_read[1]);
wire tmp_27_2;
assign tmp_27_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]);
wire tmp_27_3;
assign tmp_27_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_27_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_27_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_27_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_27_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_27_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_27_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_27_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_27_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_27_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_27_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_27_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_27_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_27_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_27_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_27_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_27_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_27_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_27_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_27_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_27_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_27_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_27_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_27_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_27_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_27_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_27_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_27_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_27_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_27_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_27_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_27_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_27_V_read[3]);
wire tmp_27_4;
assign tmp_27_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_27_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_27_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_27_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_27_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_27_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_27_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_27_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_27_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_27_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_27_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_27_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_27_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_27_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_27_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_27_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_27_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_27_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_27_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_27_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_27_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_27_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_27_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_27_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_27_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_27_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_27_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_27_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_27_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_27_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_27_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_27_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_27_V_read[4]);
wire tmp_27_5;
assign tmp_27_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]);
wire tmp_27_6;
assign tmp_27_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_27_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_27_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_27_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_27_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_27_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_27_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_27_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_27_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_27_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_27_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_27_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_27_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_27_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_27_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_27_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_27_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_27_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_27_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_27_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_27_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_27_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_27_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_27_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_27_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_27_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_27_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_27_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_27_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_27_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_27_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_27_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_27_V_read[6]);
wire tmp_27_7;
assign tmp_27_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]);
wire tmp_27_8;
assign tmp_27_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_27_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_27_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_27_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_27_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_27_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_27_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_27_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_27_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_27_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_27_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_27_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_27_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_27_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_27_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_27_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_27_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_27_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_27_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_27_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_27_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_27_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_27_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_27_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_27_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_27_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_27_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_27_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_27_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_27_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_27_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_27_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_27_V_read[8]);
wire tmp_27_9;
assign tmp_27_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_27_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_27_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_27_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_27_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_27_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_27_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_27_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_27_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_27_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_27_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_27_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_27_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_27_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_27_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_27_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_27_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_27_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_27_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_27_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_27_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_27_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_27_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_27_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_27_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_27_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_27_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_27_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_27_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_27_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_27_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_27_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_27_V_read[9]);
wire tmp_27_10;
assign tmp_27_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_27_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_27_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_27_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_27_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_27_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_27_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_27_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_27_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_27_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_27_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_27_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_27_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_27_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_27_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_27_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_27_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_27_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_27_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_27_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_27_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_27_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_27_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_27_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_27_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_27_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_27_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_27_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_27_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_27_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_27_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_27_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_27_V_read[10]);
wire tmp_27_11;
assign tmp_27_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_27_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_27_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_27_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_27_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_27_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_27_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_27_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_27_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_27_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_27_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_27_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_27_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_27_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_27_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_27_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_27_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_27_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_27_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_27_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_27_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_27_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_27_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_27_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_27_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_27_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_27_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_27_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_27_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_27_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_27_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_27_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_27_V_read[11]);
wire tmp_27_12;
assign tmp_27_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_27_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_27_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_27_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_27_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_27_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_27_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_27_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_27_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_27_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_27_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_27_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_27_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_27_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_27_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_27_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_27_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_27_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_27_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_27_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_27_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_27_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_27_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_27_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_27_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_27_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_27_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_27_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_27_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_27_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_27_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_27_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_27_V_read[12]);
wire tmp_27_13;
assign tmp_27_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_27_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_27_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_27_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_27_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_27_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_27_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_27_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_27_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_27_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_27_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_27_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_27_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_27_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_27_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_27_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_27_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_27_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_27_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_27_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_27_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_27_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_27_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_27_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_27_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_27_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_27_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_27_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_27_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_27_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_27_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_27_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_27_V_read[13]);
wire tmp_27_14;
assign tmp_27_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]);
wire tmp_27_16;
assign tmp_27_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]);
wire tmp_27_17;
assign tmp_27_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_27_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_27_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_27_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_27_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_27_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_27_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_27_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_27_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_27_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_27_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_27_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_27_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_27_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_27_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_27_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_27_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_27_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_27_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_27_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_27_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_27_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_27_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_27_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_27_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_27_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_27_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_27_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_27_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_27_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_27_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_27_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_27_V_read[17]);
wire tmp_27_18;
assign tmp_27_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_27_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_27_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_27_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_27_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_27_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_27_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_27_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_27_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_27_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_27_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_27_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_27_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_27_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_27_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_27_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_27_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_27_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_27_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_27_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_27_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_27_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_27_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_27_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_27_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_27_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_27_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_27_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_27_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_27_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_27_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_27_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_27_V_read[18]);
wire tmp_27_19;
assign tmp_27_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_27_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_27_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_27_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_27_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_27_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_27_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_27_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_27_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_27_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_27_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_27_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_27_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_27_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_27_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_27_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_27_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_27_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_27_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_27_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_27_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_27_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_27_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_27_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_27_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_27_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_27_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_27_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_27_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_27_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_27_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_27_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_27_V_read[19]);
wire tmp_27_20;
assign tmp_27_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_27_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_27_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_27_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_27_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_27_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_27_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_27_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_27_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_27_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_27_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_27_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_27_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_27_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_27_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_27_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_27_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_27_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_27_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_27_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_27_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_27_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_27_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_27_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_27_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_27_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_27_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_27_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_27_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_27_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_27_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_27_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_27_V_read[20]);
wire tmp_27_21;
assign tmp_27_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]);
wire tmp_27_22;
assign tmp_27_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_27_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_27_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_27_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_27_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_27_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_27_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_27_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_27_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_27_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_27_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_27_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_27_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_27_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_27_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_27_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_27_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_27_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_27_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_27_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_27_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_27_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_27_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_27_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_27_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_27_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_27_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_27_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_27_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_27_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_27_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_27_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_27_V_read[22]);
wire tmp_27_23;
assign tmp_27_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_27_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_27_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_27_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_27_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_27_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_27_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_27_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_27_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_27_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_27_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_27_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_27_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_27_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_27_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_27_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_27_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_27_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_27_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_27_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_27_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_27_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_27_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_27_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_27_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_27_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_27_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_27_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_27_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_27_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_27_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_27_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_27_V_read[23]);
wire tmp_27_24;
assign tmp_27_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_27_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_27_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_27_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_27_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_27_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_27_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_27_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_27_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_27_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_27_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_27_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_27_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_27_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_27_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_27_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_27_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_27_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_27_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_27_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_27_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_27_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_27_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_27_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_27_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_27_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_27_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_27_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_27_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_27_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_27_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_27_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_27_V_read[24]);
wire tmp_27_25;
assign tmp_27_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]);
wire tmp_27_26;
assign tmp_27_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_27_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_27_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_27_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_27_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_27_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_27_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_27_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_27_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_27_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_27_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_27_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_27_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_27_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_27_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_27_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_27_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_27_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_27_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_27_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_27_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_27_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_27_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_27_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_27_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_27_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_27_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_27_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_27_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_27_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_27_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_27_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_27_V_read[26]);
wire tmp_27_27;
assign tmp_27_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_27_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_27_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_27_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_27_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_27_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_27_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_27_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_27_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_27_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_27_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_27_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_27_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_27_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_27_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_27_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_27_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_27_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_27_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_27_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_27_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_27_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_27_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_27_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_27_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_27_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_27_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_27_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_27_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_27_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_27_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_27_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_27_V_read[27]);
wire tmp_27_29;
assign tmp_27_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_27_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_27_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_27_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_27_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_27_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_27_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_27_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_27_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_27_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_27_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_27_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_27_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_27_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_27_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_27_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_27_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_27_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_27_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_27_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_27_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_27_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_27_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_27_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_27_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_27_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_27_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_27_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_27_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_27_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_27_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_27_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_27_V_read[29]);
wire tmp_27_30;
assign tmp_27_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_27_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_27_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_27_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_27_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_27_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_27_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_27_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_27_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_27_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_27_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_27_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_27_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_27_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_27_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_27_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_27_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_27_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_27_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_27_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_27_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_27_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_27_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_27_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_27_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_27_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_27_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_27_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_27_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_27_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_27_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_27_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_27_V_read[30]);
wire tmp_27_31;
assign tmp_27_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]);
assign ap_return_27 = {tmp_27_0,tmp_27_1,tmp_27_2,tmp_27_3,tmp_27_4,tmp_27_5,tmp_27_6,tmp_27_7,tmp_27_8,tmp_27_9,tmp_27_10,tmp_27_11,tmp_27_12,tmp_27_13,tmp_27_14,1'b0,tmp_27_16,tmp_27_17,tmp_27_18,tmp_27_19,tmp_27_20,tmp_27_21,tmp_27_22,tmp_27_23,tmp_27_24,tmp_27_25,tmp_27_26,tmp_27_27,1'b0,tmp_27_29,tmp_27_30,tmp_27_31};
wire tmp_28_0;
assign tmp_28_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]);
wire tmp_28_1;
assign tmp_28_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_28_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_28_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_28_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_28_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_28_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_28_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_28_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_28_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_28_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_28_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_28_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_28_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_28_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_28_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_28_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_28_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_28_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_28_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_28_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_28_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_28_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_28_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_28_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_28_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_28_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_28_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_28_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_28_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_28_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_28_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_28_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_28_V_read[1]);
wire tmp_28_2;
assign tmp_28_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_28_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_28_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_28_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_28_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_28_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_28_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_28_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_28_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_28_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_28_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_28_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_28_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_28_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_28_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_28_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_28_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_28_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_28_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_28_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_28_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_28_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_28_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_28_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_28_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_28_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_28_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_28_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_28_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_28_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_28_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_28_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_28_V_read[2]);
wire tmp_28_3;
assign tmp_28_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]);
wire tmp_28_5;
assign tmp_28_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_28_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_28_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_28_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_28_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_28_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_28_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_28_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_28_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_28_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_28_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_28_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_28_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_28_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_28_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_28_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_28_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_28_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_28_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_28_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_28_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_28_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_28_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_28_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_28_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_28_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_28_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_28_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_28_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_28_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_28_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_28_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_28_V_read[5]);
wire tmp_28_6;
assign tmp_28_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_28_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_28_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_28_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_28_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_28_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_28_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_28_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_28_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_28_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_28_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_28_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_28_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_28_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_28_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_28_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_28_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_28_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_28_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_28_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_28_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_28_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_28_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_28_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_28_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_28_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_28_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_28_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_28_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_28_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_28_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_28_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_28_V_read[6]);
wire tmp_28_7;
assign tmp_28_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]);
wire tmp_28_8;
assign tmp_28_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_28_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_28_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_28_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_28_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_28_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_28_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_28_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_28_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_28_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_28_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_28_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_28_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_28_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_28_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_28_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_28_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_28_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_28_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_28_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_28_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_28_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_28_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_28_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_28_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_28_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_28_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_28_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_28_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_28_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_28_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_28_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_28_V_read[8]);
wire tmp_28_9;
assign tmp_28_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_28_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_28_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_28_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_28_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_28_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_28_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_28_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_28_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_28_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_28_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_28_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_28_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_28_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_28_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_28_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_28_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_28_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_28_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_28_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_28_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_28_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_28_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_28_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_28_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_28_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_28_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_28_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_28_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_28_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_28_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_28_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_28_V_read[9]);
wire tmp_28_10;
assign tmp_28_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_28_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_28_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_28_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_28_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_28_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_28_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_28_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_28_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_28_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_28_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_28_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_28_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_28_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_28_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_28_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_28_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_28_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_28_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_28_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_28_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_28_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_28_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_28_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_28_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_28_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_28_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_28_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_28_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_28_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_28_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_28_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_28_V_read[10]);
wire tmp_28_11;
assign tmp_28_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_28_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_28_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_28_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_28_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_28_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_28_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_28_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_28_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_28_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_28_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_28_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_28_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_28_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_28_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_28_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_28_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_28_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_28_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_28_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_28_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_28_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_28_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_28_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_28_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_28_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_28_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_28_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_28_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_28_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_28_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_28_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_28_V_read[11]);
wire tmp_28_12;
assign tmp_28_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_28_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_28_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_28_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_28_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_28_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_28_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_28_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_28_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_28_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_28_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_28_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_28_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_28_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_28_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_28_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_28_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_28_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_28_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_28_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_28_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_28_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_28_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_28_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_28_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_28_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_28_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_28_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_28_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_28_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_28_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_28_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_28_V_read[12]);
wire tmp_28_13;
assign tmp_28_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]);
wire tmp_28_14;
assign tmp_28_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_28_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_28_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_28_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_28_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_28_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_28_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_28_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_28_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_28_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_28_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_28_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_28_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_28_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_28_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_28_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_28_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_28_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_28_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_28_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_28_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_28_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_28_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_28_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_28_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_28_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_28_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_28_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_28_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_28_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_28_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_28_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_28_V_read[14]);
wire tmp_28_16;
assign tmp_28_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]);
wire tmp_28_17;
assign tmp_28_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_28_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_28_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_28_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_28_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_28_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_28_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_28_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_28_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_28_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_28_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_28_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_28_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_28_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_28_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_28_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_28_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_28_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_28_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_28_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_28_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_28_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_28_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_28_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_28_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_28_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_28_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_28_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_28_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_28_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_28_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_28_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_28_V_read[17]);
wire tmp_28_18;
assign tmp_28_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_28_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_28_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_28_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_28_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_28_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_28_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_28_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_28_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_28_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_28_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_28_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_28_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_28_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_28_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_28_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_28_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_28_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_28_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_28_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_28_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_28_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_28_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_28_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_28_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_28_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_28_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_28_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_28_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_28_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_28_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_28_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_28_V_read[18]);
wire tmp_28_19;
assign tmp_28_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_28_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_28_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_28_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_28_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_28_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_28_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_28_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_28_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_28_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_28_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_28_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_28_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_28_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_28_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_28_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_28_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_28_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_28_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_28_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_28_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_28_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_28_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_28_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_28_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_28_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_28_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_28_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_28_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_28_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_28_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_28_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_28_V_read[19]);
wire tmp_28_20;
assign tmp_28_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_28_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_28_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_28_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_28_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_28_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_28_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_28_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_28_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_28_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_28_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_28_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_28_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_28_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_28_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_28_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_28_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_28_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_28_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_28_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_28_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_28_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_28_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_28_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_28_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_28_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_28_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_28_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_28_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_28_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_28_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_28_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_28_V_read[20]);
wire tmp_28_21;
assign tmp_28_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]);
wire tmp_28_23;
assign tmp_28_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_28_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_28_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_28_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_28_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_28_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_28_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_28_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_28_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_28_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_28_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_28_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_28_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_28_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_28_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_28_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_28_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_28_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_28_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_28_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_28_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_28_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_28_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_28_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_28_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_28_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_28_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_28_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_28_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_28_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_28_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_28_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_28_V_read[23]);
wire tmp_28_24;
assign tmp_28_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]);
wire tmp_28_25;
assign tmp_28_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_28_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_28_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_28_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_28_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_28_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_28_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_28_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_28_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_28_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_28_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_28_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_28_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_28_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_28_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_28_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_28_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_28_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_28_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_28_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_28_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_28_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_28_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_28_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_28_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_28_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_28_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_28_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_28_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_28_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_28_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_28_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_28_V_read[25]);
wire tmp_28_26;
assign tmp_28_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]);
wire tmp_28_27;
assign tmp_28_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_28_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_28_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_28_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_28_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_28_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_28_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_28_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_28_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_28_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_28_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_28_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_28_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_28_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_28_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_28_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_28_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_28_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_28_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_28_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_28_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_28_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_28_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_28_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_28_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_28_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_28_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_28_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_28_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_28_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_28_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_28_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_28_V_read[27]);
wire tmp_28_28;
assign tmp_28_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]);
wire tmp_28_30;
assign tmp_28_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]);
wire tmp_28_31;
assign tmp_28_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]);
assign ap_return_28 = {tmp_28_0,tmp_28_1,tmp_28_2,tmp_28_3,1'b0,tmp_28_5,tmp_28_6,tmp_28_7,tmp_28_8,tmp_28_9,tmp_28_10,tmp_28_11,tmp_28_12,tmp_28_13,tmp_28_14,1'b0,tmp_28_16,tmp_28_17,tmp_28_18,tmp_28_19,tmp_28_20,tmp_28_21,1'b0,tmp_28_23,tmp_28_24,tmp_28_25,tmp_28_26,tmp_28_27,tmp_28_28,1'b0,tmp_28_30,tmp_28_31};
wire tmp_29_0;
assign tmp_29_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]);
wire tmp_29_1;
assign tmp_29_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_29_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_29_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_29_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_29_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_29_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_29_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_29_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_29_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_29_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_29_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_29_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_29_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_29_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_29_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_29_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_29_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_29_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_29_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_29_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_29_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_29_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_29_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_29_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_29_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_29_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_29_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_29_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_29_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_29_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_29_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_29_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_29_V_read[1]);
wire tmp_29_2;
assign tmp_29_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_29_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_29_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_29_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_29_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_29_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_29_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_29_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_29_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_29_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_29_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_29_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_29_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_29_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_29_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_29_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_29_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_29_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_29_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_29_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_29_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_29_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_29_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_29_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_29_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_29_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_29_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_29_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_29_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_29_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_29_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_29_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_29_V_read[2]);
wire tmp_29_3;
assign tmp_29_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_29_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_29_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_29_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_29_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_29_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_29_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_29_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_29_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_29_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_29_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_29_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_29_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_29_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_29_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_29_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_29_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_29_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_29_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_29_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_29_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_29_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_29_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_29_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_29_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_29_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_29_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_29_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_29_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_29_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_29_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_29_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_29_V_read[3]);
wire tmp_29_4;
assign tmp_29_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_29_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_29_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_29_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_29_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_29_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_29_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_29_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_29_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_29_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_29_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_29_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_29_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_29_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_29_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_29_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_29_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_29_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_29_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_29_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_29_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_29_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_29_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_29_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_29_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_29_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_29_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_29_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_29_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_29_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_29_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_29_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_29_V_read[4]);
wire tmp_29_5;
assign tmp_29_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_29_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_29_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_29_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_29_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_29_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_29_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_29_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_29_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_29_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_29_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_29_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_29_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_29_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_29_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_29_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_29_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_29_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_29_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_29_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_29_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_29_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_29_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_29_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_29_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_29_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_29_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_29_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_29_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_29_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_29_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_29_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_29_V_read[5]);
wire tmp_29_6;
assign tmp_29_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_29_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_29_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_29_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_29_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_29_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_29_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_29_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_29_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_29_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_29_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_29_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_29_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_29_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_29_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_29_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_29_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_29_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_29_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_29_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_29_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_29_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_29_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_29_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_29_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_29_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_29_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_29_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_29_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_29_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_29_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_29_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_29_V_read[6]);
wire tmp_29_7;
assign tmp_29_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]);
wire tmp_29_8;
assign tmp_29_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_29_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_29_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_29_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_29_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_29_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_29_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_29_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_29_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_29_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_29_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_29_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_29_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_29_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_29_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_29_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_29_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_29_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_29_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_29_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_29_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_29_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_29_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_29_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_29_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_29_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_29_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_29_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_29_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_29_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_29_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_29_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_29_V_read[8]);
wire tmp_29_9;
assign tmp_29_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_29_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_29_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_29_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_29_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_29_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_29_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_29_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_29_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_29_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_29_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_29_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_29_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_29_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_29_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_29_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_29_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_29_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_29_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_29_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_29_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_29_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_29_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_29_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_29_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_29_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_29_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_29_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_29_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_29_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_29_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_29_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_29_V_read[9]);
wire tmp_29_10;
assign tmp_29_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_29_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_29_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_29_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_29_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_29_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_29_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_29_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_29_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_29_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_29_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_29_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_29_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_29_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_29_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_29_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_29_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_29_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_29_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_29_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_29_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_29_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_29_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_29_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_29_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_29_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_29_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_29_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_29_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_29_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_29_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_29_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_29_V_read[10]);
wire tmp_29_11;
assign tmp_29_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]);
wire tmp_29_12;
assign tmp_29_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_29_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_29_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_29_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_29_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_29_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_29_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_29_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_29_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_29_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_29_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_29_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_29_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_29_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_29_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_29_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_29_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_29_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_29_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_29_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_29_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_29_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_29_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_29_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_29_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_29_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_29_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_29_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_29_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_29_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_29_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_29_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_29_V_read[12]);
wire tmp_29_13;
assign tmp_29_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_29_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_29_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_29_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_29_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_29_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_29_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_29_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_29_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_29_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_29_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_29_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_29_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_29_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_29_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_29_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_29_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_29_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_29_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_29_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_29_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_29_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_29_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_29_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_29_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_29_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_29_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_29_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_29_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_29_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_29_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_29_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_29_V_read[13]);
wire tmp_29_14;
assign tmp_29_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_29_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_29_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_29_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_29_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_29_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_29_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_29_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_29_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_29_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_29_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_29_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_29_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_29_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_29_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_29_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_29_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_29_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_29_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_29_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_29_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_29_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_29_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_29_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_29_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_29_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_29_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_29_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_29_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_29_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_29_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_29_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_29_V_read[14]);
wire tmp_29_15;
assign tmp_29_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_29_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_29_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_29_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_29_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_29_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_29_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_29_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_29_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_29_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_29_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_29_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_29_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_29_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_29_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_29_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_29_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_29_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_29_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_29_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_29_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_29_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_29_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_29_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_29_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_29_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_29_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_29_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_29_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_29_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_29_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_29_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_29_V_read[15]);
wire tmp_29_16;
assign tmp_29_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]);
wire tmp_29_17;
assign tmp_29_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]);
wire tmp_29_18;
assign tmp_29_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_29_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_29_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_29_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_29_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_29_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_29_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_29_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_29_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_29_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_29_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_29_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_29_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_29_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_29_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_29_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_29_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_29_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_29_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_29_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_29_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_29_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_29_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_29_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_29_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_29_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_29_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_29_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_29_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_29_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_29_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_29_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_29_V_read[18]);
wire tmp_29_19;
assign tmp_29_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_29_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_29_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_29_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_29_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_29_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_29_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_29_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_29_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_29_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_29_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_29_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_29_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_29_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_29_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_29_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_29_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_29_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_29_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_29_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_29_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_29_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_29_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_29_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_29_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_29_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_29_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_29_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_29_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_29_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_29_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_29_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_29_V_read[19]);
wire tmp_29_20;
assign tmp_29_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_29_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_29_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_29_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_29_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_29_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_29_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_29_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_29_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_29_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_29_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_29_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_29_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_29_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_29_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_29_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_29_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_29_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_29_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_29_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_29_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_29_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_29_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_29_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_29_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_29_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_29_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_29_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_29_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_29_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_29_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_29_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_29_V_read[20]);
wire tmp_29_21;
assign tmp_29_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_29_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_29_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_29_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_29_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_29_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_29_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_29_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_29_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_29_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_29_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_29_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_29_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_29_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_29_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_29_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_29_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_29_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_29_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_29_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_29_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_29_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_29_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_29_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_29_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_29_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_29_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_29_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_29_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_29_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_29_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_29_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_29_V_read[21]);
wire tmp_29_22;
assign tmp_29_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]);
wire tmp_29_23;
assign tmp_29_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]);
wire tmp_29_24;
assign tmp_29_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_29_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_29_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_29_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_29_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_29_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_29_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_29_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_29_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_29_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_29_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_29_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_29_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_29_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_29_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_29_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_29_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_29_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_29_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_29_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_29_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_29_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_29_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_29_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_29_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_29_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_29_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_29_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_29_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_29_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_29_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_29_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_29_V_read[24]);
wire tmp_29_25;
assign tmp_29_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]);
wire tmp_29_26;
assign tmp_29_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_29_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_29_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_29_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_29_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_29_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_29_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_29_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_29_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_29_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_29_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_29_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_29_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_29_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_29_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_29_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_29_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_29_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_29_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_29_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_29_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_29_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_29_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_29_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_29_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_29_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_29_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_29_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_29_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_29_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_29_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_29_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_29_V_read[26]);
wire tmp_29_27;
assign tmp_29_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_29_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_29_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_29_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_29_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_29_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_29_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_29_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_29_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_29_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_29_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_29_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_29_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_29_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_29_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_29_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_29_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_29_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_29_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_29_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_29_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_29_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_29_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_29_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_29_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_29_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_29_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_29_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_29_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_29_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_29_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_29_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_29_V_read[27]);
wire tmp_29_28;
assign tmp_29_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_29_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_29_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_29_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_29_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_29_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_29_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_29_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_29_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_29_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_29_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_29_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_29_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_29_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_29_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_29_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_29_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_29_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_29_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_29_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_29_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_29_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_29_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_29_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_29_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_29_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_29_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_29_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_29_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_29_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_29_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_29_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_29_V_read[28]);
wire tmp_29_29;
assign tmp_29_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]);
wire tmp_29_31;
assign tmp_29_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_29_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_29_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_29_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_29_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_29_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_29_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_29_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_29_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_29_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_29_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_29_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_29_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_29_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_29_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_29_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_29_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_29_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_29_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_29_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_29_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_29_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_29_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_29_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_29_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_29_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_29_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_29_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_29_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_29_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_29_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_29_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_29_V_read[31]);
assign ap_return_29 = {tmp_29_0,tmp_29_1,tmp_29_2,tmp_29_3,tmp_29_4,tmp_29_5,tmp_29_6,tmp_29_7,tmp_29_8,tmp_29_9,tmp_29_10,tmp_29_11,tmp_29_12,tmp_29_13,tmp_29_14,tmp_29_15,tmp_29_16,tmp_29_17,tmp_29_18,tmp_29_19,tmp_29_20,tmp_29_21,tmp_29_22,tmp_29_23,tmp_29_24,tmp_29_25,tmp_29_26,tmp_29_27,tmp_29_28,tmp_29_29,1'b0,tmp_29_31};
wire tmp_30_0;
assign tmp_30_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]);
wire tmp_30_1;
assign tmp_30_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_30_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_30_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_30_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_30_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_30_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_30_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_30_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_30_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_30_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_30_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_30_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_30_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_30_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_30_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_30_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_30_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_30_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_30_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_30_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_30_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_30_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_30_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_30_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_30_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_30_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_30_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_30_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_30_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_30_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_30_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_30_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_30_V_read[1]);
wire tmp_30_2;
assign tmp_30_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_30_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_30_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_30_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_30_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_30_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_30_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_30_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_30_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_30_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_30_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_30_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_30_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_30_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_30_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_30_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_30_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_30_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_30_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_30_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_30_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_30_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_30_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_30_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_30_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_30_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_30_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_30_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_30_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_30_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_30_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_30_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_30_V_read[2]);
wire tmp_30_3;
assign tmp_30_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]);
wire tmp_30_4;
assign tmp_30_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_30_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_30_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_30_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_30_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_30_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_30_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_30_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_30_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_30_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_30_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_30_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_30_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_30_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_30_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_30_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_30_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_30_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_30_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_30_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_30_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_30_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_30_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_30_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_30_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_30_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_30_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_30_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_30_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_30_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_30_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_30_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_30_V_read[4]);
wire tmp_30_5;
assign tmp_30_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_30_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_30_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_30_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_30_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_30_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_30_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_30_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_30_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_30_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_30_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_30_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_30_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_30_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_30_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_30_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_30_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_30_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_30_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_30_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_30_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_30_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_30_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_30_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_30_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_30_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_30_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_30_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_30_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_30_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_30_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_30_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_30_V_read[5]);
wire tmp_30_6;
assign tmp_30_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]);
wire tmp_30_7;
assign tmp_30_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_30_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_30_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_30_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_30_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_30_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_30_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_30_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_30_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_30_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_30_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_30_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_30_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_30_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_30_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_30_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_30_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_30_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_30_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_30_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_30_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_30_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_30_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_30_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_30_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_30_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_30_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_30_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_30_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_30_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_30_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_30_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_30_V_read[7]);
wire tmp_30_8;
assign tmp_30_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]);
wire tmp_30_9;
assign tmp_30_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]);
wire tmp_30_10;
assign tmp_30_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]);
wire tmp_30_11;
assign tmp_30_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]);
wire tmp_30_13;
assign tmp_30_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_30_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_30_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_30_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_30_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_30_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_30_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_30_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_30_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_30_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_30_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_30_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_30_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_30_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_30_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_30_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_30_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_30_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_30_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_30_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_30_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_30_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_30_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_30_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_30_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_30_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_30_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_30_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_30_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_30_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_30_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_30_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_30_V_read[13]);
wire tmp_30_14;
assign tmp_30_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_30_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_30_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_30_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_30_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_30_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_30_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_30_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_30_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_30_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_30_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_30_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_30_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_30_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_30_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_30_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_30_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_30_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_30_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_30_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_30_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_30_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_30_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_30_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_30_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_30_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_30_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_30_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_30_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_30_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_30_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_30_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_30_V_read[14]);
wire tmp_30_15;
assign tmp_30_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_30_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_30_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_30_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_30_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_30_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_30_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_30_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_30_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_30_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_30_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_30_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_30_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_30_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_30_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_30_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_30_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_30_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_30_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_30_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_30_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_30_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_30_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_30_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_30_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_30_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_30_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_30_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_30_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_30_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_30_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_30_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_30_V_read[15]);
wire tmp_30_16;
assign tmp_30_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_30_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_30_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_30_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_30_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_30_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_30_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_30_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_30_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_30_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_30_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_30_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_30_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_30_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_30_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_30_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_30_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_30_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_30_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_30_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_30_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_30_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_30_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_30_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_30_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_30_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_30_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_30_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_30_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_30_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_30_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_30_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_30_V_read[16]);
wire tmp_30_18;
assign tmp_30_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_30_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_30_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_30_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_30_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_30_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_30_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_30_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_30_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_30_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_30_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_30_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_30_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_30_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_30_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_30_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_30_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_30_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_30_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_30_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_30_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_30_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_30_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_30_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_30_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_30_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_30_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_30_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_30_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_30_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_30_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_30_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_30_V_read[18]);
wire tmp_30_19;
assign tmp_30_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]);
wire tmp_30_20;
assign tmp_30_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_30_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_30_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_30_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_30_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_30_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_30_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_30_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_30_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_30_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_30_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_30_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_30_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_30_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_30_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_30_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_30_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_30_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_30_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_30_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_30_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_30_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_30_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_30_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_30_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_30_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_30_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_30_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_30_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_30_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_30_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_30_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_30_V_read[20]);
wire tmp_30_21;
assign tmp_30_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]);
wire tmp_30_22;
assign tmp_30_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_30_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_30_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_30_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_30_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_30_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_30_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_30_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_30_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_30_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_30_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_30_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_30_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_30_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_30_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_30_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_30_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_30_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_30_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_30_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_30_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_30_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_30_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_30_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_30_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_30_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_30_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_30_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_30_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_30_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_30_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_30_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_30_V_read[22]);
wire tmp_30_23;
assign tmp_30_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_30_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_30_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_30_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_30_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_30_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_30_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_30_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_30_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_30_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_30_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_30_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_30_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_30_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_30_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_30_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_30_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_30_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_30_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_30_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_30_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_30_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_30_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_30_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_30_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_30_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_30_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_30_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_30_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_30_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_30_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_30_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_30_V_read[23]);
wire tmp_30_24;
assign tmp_30_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]);
wire tmp_30_25;
assign tmp_30_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]);
wire tmp_30_26;
assign tmp_30_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_30_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_30_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_30_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_30_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_30_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_30_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_30_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_30_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_30_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_30_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_30_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_30_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_30_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_30_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_30_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_30_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_30_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_30_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_30_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_30_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_30_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_30_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_30_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_30_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_30_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_30_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_30_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_30_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_30_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_30_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_30_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_30_V_read[26]);
wire tmp_30_27;
assign tmp_30_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_30_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_30_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_30_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_30_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_30_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_30_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_30_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_30_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_30_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_30_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_30_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_30_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_30_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_30_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_30_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_30_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_30_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_30_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_30_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_30_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_30_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_30_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_30_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_30_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_30_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_30_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_30_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_30_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_30_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_30_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_30_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_30_V_read[27]);
wire tmp_30_28;
assign tmp_30_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_30_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_30_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_30_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_30_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_30_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_30_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_30_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_30_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_30_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_30_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_30_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_30_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_30_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_30_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_30_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_30_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_30_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_30_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_30_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_30_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_30_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_30_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_30_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_30_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_30_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_30_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_30_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_30_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_30_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_30_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_30_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_30_V_read[28]);
wire tmp_30_29;
assign tmp_30_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_30_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_30_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_30_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_30_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_30_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_30_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_30_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_30_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_30_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_30_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_30_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_30_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_30_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_30_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_30_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_30_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_30_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_30_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_30_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_30_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_30_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_30_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_30_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_30_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_30_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_30_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_30_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_30_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_30_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_30_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_30_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_30_V_read[29]);
wire tmp_30_31;
assign tmp_30_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]);
assign ap_return_30 = {tmp_30_0,tmp_30_1,tmp_30_2,tmp_30_3,tmp_30_4,tmp_30_5,tmp_30_6,tmp_30_7,tmp_30_8,tmp_30_9,tmp_30_10,tmp_30_11,1'b0,tmp_30_13,tmp_30_14,tmp_30_15,tmp_30_16,1'b0,tmp_30_18,tmp_30_19,tmp_30_20,tmp_30_21,tmp_30_22,tmp_30_23,tmp_30_24,tmp_30_25,tmp_30_26,tmp_30_27,tmp_30_28,tmp_30_29,1'b0,tmp_30_31};
wire tmp_31_0;
assign tmp_31_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]);
wire tmp_31_1;
assign tmp_31_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_31_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_31_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_31_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_31_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_31_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_31_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_31_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_31_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_31_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_31_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_31_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_31_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_31_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_31_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_31_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_31_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_31_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_31_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_31_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_31_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_31_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_31_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_31_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_31_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_31_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_31_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_31_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_31_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_31_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_31_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_31_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_31_V_read[1]);
wire tmp_31_2;
assign tmp_31_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_31_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_31_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_31_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_31_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_31_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_31_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_31_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_31_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_31_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_31_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_31_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_31_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_31_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_31_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_31_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_31_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_31_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_31_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_31_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_31_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_31_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_31_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_31_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_31_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_31_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_31_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_31_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_31_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_31_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_31_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_31_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_31_V_read[2]);
wire tmp_31_3;
assign tmp_31_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]);
wire tmp_31_4;
assign tmp_31_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_31_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_31_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_31_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_31_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_31_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_31_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_31_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_31_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_31_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_31_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_31_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_31_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_31_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_31_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_31_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_31_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_31_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_31_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_31_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_31_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_31_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_31_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_31_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_31_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_31_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_31_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_31_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_31_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_31_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_31_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_31_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_31_V_read[4]);
wire tmp_31_5;
assign tmp_31_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_31_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_31_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_31_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_31_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_31_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_31_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_31_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_31_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_31_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_31_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_31_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_31_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_31_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_31_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_31_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_31_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_31_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_31_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_31_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_31_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_31_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_31_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_31_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_31_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_31_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_31_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_31_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_31_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_31_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_31_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_31_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_31_V_read[5]);
wire tmp_31_6;
assign tmp_31_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_31_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_31_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_31_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_31_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_31_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_31_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_31_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_31_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_31_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_31_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_31_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_31_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_31_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_31_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_31_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_31_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_31_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_31_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_31_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_31_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_31_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_31_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_31_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_31_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_31_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_31_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_31_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_31_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_31_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_31_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_31_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_31_V_read[6]);
wire tmp_31_7;
assign tmp_31_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]);
wire tmp_31_8;
assign tmp_31_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]);
wire tmp_31_9;
assign tmp_31_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_31_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_31_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_31_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_31_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_31_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_31_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_31_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_31_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_31_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_31_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_31_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_31_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_31_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_31_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_31_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_31_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_31_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_31_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_31_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_31_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_31_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_31_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_31_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_31_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_31_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_31_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_31_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_31_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_31_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_31_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_31_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_31_V_read[9]);
wire tmp_31_11;
assign tmp_31_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_31_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_31_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_31_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_31_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_31_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_31_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_31_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_31_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_31_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_31_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_31_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_31_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_31_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_31_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_31_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_31_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_31_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_31_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_31_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_31_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_31_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_31_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_31_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_31_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_31_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_31_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_31_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_31_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_31_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_31_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_31_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_31_V_read[11]);
wire tmp_31_12;
assign tmp_31_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_31_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_31_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_31_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_31_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_31_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_31_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_31_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_31_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_31_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_31_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_31_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_31_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_31_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_31_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_31_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_31_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_31_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_31_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_31_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_31_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_31_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_31_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_31_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_31_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_31_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_31_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_31_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_31_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_31_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_31_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_31_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_31_V_read[12]);
wire tmp_31_13;
assign tmp_31_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_31_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_31_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_31_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_31_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_31_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_31_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_31_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_31_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_31_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_31_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_31_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_31_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_31_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_31_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_31_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_31_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_31_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_31_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_31_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_31_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_31_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_31_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_31_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_31_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_31_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_31_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_31_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_31_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_31_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_31_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_31_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_31_V_read[13]);
wire tmp_31_14;
assign tmp_31_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_31_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_31_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_31_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_31_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_31_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_31_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_31_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_31_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_31_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_31_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_31_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_31_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_31_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_31_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_31_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_31_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_31_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_31_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_31_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_31_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_31_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_31_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_31_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_31_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_31_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_31_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_31_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_31_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_31_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_31_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_31_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_31_V_read[14]);
wire tmp_31_16;
assign tmp_31_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_31_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_31_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_31_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_31_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_31_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_31_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_31_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_31_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_31_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_31_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_31_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_31_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_31_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_31_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_31_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_31_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_31_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_31_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_31_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_31_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_31_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_31_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_31_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_31_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_31_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_31_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_31_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_31_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_31_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_31_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_31_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_31_V_read[16]);
wire tmp_31_17;
assign tmp_31_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_31_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_31_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_31_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_31_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_31_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_31_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_31_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_31_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_31_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_31_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_31_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_31_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_31_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_31_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_31_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_31_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_31_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_31_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_31_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_31_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_31_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_31_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_31_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_31_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_31_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_31_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_31_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_31_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_31_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_31_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_31_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_31_V_read[17]);
wire tmp_31_18;
assign tmp_31_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_31_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_31_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_31_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_31_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_31_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_31_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_31_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_31_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_31_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_31_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_31_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_31_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_31_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_31_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_31_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_31_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_31_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_31_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_31_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_31_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_31_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_31_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_31_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_31_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_31_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_31_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_31_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_31_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_31_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_31_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_31_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_31_V_read[18]);
wire tmp_31_19;
assign tmp_31_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_31_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_31_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_31_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_31_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_31_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_31_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_31_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_31_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_31_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_31_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_31_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_31_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_31_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_31_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_31_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_31_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_31_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_31_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_31_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_31_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_31_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_31_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_31_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_31_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_31_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_31_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_31_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_31_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_31_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_31_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_31_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_31_V_read[19]);
wire tmp_31_20;
assign tmp_31_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_31_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_31_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_31_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_31_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_31_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_31_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_31_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_31_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_31_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_31_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_31_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_31_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_31_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_31_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_31_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_31_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_31_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_31_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_31_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_31_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_31_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_31_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_31_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_31_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_31_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_31_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_31_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_31_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_31_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_31_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_31_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_31_V_read[20]);
wire tmp_31_21;
assign tmp_31_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_31_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_31_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_31_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_31_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_31_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_31_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_31_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_31_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_31_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_31_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_31_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_31_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_31_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_31_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_31_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_31_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_31_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_31_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_31_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_31_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_31_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_31_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_31_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_31_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_31_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_31_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_31_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_31_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_31_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_31_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_31_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_31_V_read[21]);
wire tmp_31_22;
assign tmp_31_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_31_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_31_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_31_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_31_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_31_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_31_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_31_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_31_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_31_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_31_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_31_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_31_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_31_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_31_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_31_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_31_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_31_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_31_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_31_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_31_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_31_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_31_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_31_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_31_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_31_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_31_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_31_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_31_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_31_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_31_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_31_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_31_V_read[22]);
wire tmp_31_23;
assign tmp_31_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]);
wire tmp_31_24;
assign tmp_31_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_31_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_31_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_31_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_31_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_31_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_31_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_31_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_31_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_31_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_31_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_31_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_31_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_31_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_31_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_31_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_31_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_31_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_31_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_31_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_31_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_31_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_31_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_31_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_31_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_31_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_31_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_31_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_31_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_31_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_31_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_31_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_31_V_read[24]);
wire tmp_31_25;
assign tmp_31_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_31_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_31_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_31_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_31_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_31_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_31_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_31_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_31_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_31_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_31_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_31_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_31_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_31_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_31_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_31_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_31_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_31_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_31_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_31_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_31_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_31_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_31_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_31_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_31_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_31_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_31_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_31_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_31_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_31_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_31_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_31_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_31_V_read[25]);
wire tmp_31_26;
assign tmp_31_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_31_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_31_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_31_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_31_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_31_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_31_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_31_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_31_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_31_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_31_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_31_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_31_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_31_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_31_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_31_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_31_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_31_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_31_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_31_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_31_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_31_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_31_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_31_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_31_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_31_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_31_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_31_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_31_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_31_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_31_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_31_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_31_V_read[26]);
wire tmp_31_27;
assign tmp_31_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_31_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_31_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_31_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_31_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_31_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_31_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_31_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_31_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_31_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_31_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_31_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_31_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_31_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_31_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_31_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_31_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_31_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_31_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_31_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_31_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_31_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_31_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_31_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_31_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_31_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_31_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_31_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_31_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_31_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_31_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_31_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_31_V_read[27]);
wire tmp_31_28;
assign tmp_31_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]);
wire tmp_31_29;
assign tmp_31_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]);
wire tmp_31_30;
assign tmp_31_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_31_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_31_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_31_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_31_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_31_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_31_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_31_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_31_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_31_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_31_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_31_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_31_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_31_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_31_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_31_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_31_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_31_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_31_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_31_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_31_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_31_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_31_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_31_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_31_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_31_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_31_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_31_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_31_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_31_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_31_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_31_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_31_V_read[30]);
wire tmp_31_31;
assign tmp_31_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]);
assign ap_return_31 = {tmp_31_0,tmp_31_1,tmp_31_2,tmp_31_3,tmp_31_4,tmp_31_5,tmp_31_6,tmp_31_7,tmp_31_8,tmp_31_9,1'b0,tmp_31_11,tmp_31_12,tmp_31_13,tmp_31_14,1'b0,tmp_31_16,tmp_31_17,tmp_31_18,tmp_31_19,tmp_31_20,tmp_31_21,tmp_31_22,tmp_31_23,tmp_31_24,tmp_31_25,tmp_31_26,tmp_31_27,tmp_31_28,tmp_31_29,tmp_31_30,tmp_31_31};
endmodule