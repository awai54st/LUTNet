`timescale 1 ns / 1 ps

module LUTARRAY (
        in_V,
        in_1_V,
        in_2_V,
        in_3_V,
        weight_0_0_V_read,
        weight_0_1_V_read,
        weight_0_2_V_read,
        weight_0_3_V_read,
        weight_0_4_V_read,
        weight_0_5_V_read,
        weight_0_6_V_read,
        weight_0_7_V_read,
        weight_0_8_V_read,
        weight_0_9_V_read,
        weight_0_10_V_read,
        weight_0_11_V_read,
        weight_0_12_V_read,
        weight_0_13_V_read,
        weight_0_14_V_read,
        weight_0_15_V_read,
        weight_0_16_V_read,
        weight_0_17_V_read,
        weight_0_18_V_read,
        weight_0_19_V_read,
        weight_0_20_V_read,
        weight_0_21_V_read,
        weight_0_22_V_read,
        weight_0_23_V_read,
        weight_0_24_V_read,
        weight_0_25_V_read,
        weight_0_26_V_read,
        weight_0_27_V_read,
        weight_0_28_V_read,
        weight_0_29_V_read,
        weight_0_30_V_read,
        weight_0_31_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15,
        ap_return_16,
        ap_return_17,
        ap_return_18,
        ap_return_19,
        ap_return_20,
        ap_return_21,
        ap_return_22,
        ap_return_23,
        ap_return_24,
        ap_return_25,
        ap_return_26,
        ap_return_27,
        ap_return_28,
        ap_return_29,
        ap_return_30,
        ap_return_31);



input  [31:0] in_V;
input  [31:0] in_1_V;
input  [31:0] in_2_V;
input  [31:0] in_3_V;
input  [31:0] weight_0_0_V_read;
input  [31:0] weight_0_1_V_read;
input  [31:0] weight_0_2_V_read;
input  [31:0] weight_0_3_V_read;
input  [31:0] weight_0_4_V_read;
input  [31:0] weight_0_5_V_read;
input  [31:0] weight_0_6_V_read;
input  [31:0] weight_0_7_V_read;
input  [31:0] weight_0_8_V_read;
input  [31:0] weight_0_9_V_read;
input  [31:0] weight_0_10_V_read;
input  [31:0] weight_0_11_V_read;
input  [31:0] weight_0_12_V_read;
input  [31:0] weight_0_13_V_read;
input  [31:0] weight_0_14_V_read;
input  [31:0] weight_0_15_V_read;
input  [31:0] weight_0_16_V_read;
input  [31:0] weight_0_17_V_read;
input  [31:0] weight_0_18_V_read;
input  [31:0] weight_0_19_V_read;
input  [31:0] weight_0_20_V_read;
input  [31:0] weight_0_21_V_read;
input  [31:0] weight_0_22_V_read;
input  [31:0] weight_0_23_V_read;
input  [31:0] weight_0_24_V_read;
input  [31:0] weight_0_25_V_read;
input  [31:0] weight_0_26_V_read;
input  [31:0] weight_0_27_V_read;
input  [31:0] weight_0_28_V_read;
input  [31:0] weight_0_29_V_read;
input  [31:0] weight_0_30_V_read;
input  [31:0] weight_0_31_V_read;
output  [31:0] ap_return_0;
output  [31:0] ap_return_1;
output  [31:0] ap_return_2;
output  [31:0] ap_return_3;
output  [31:0] ap_return_4;
output  [31:0] ap_return_5;
output  [31:0] ap_return_6;
output  [31:0] ap_return_7;
output  [31:0] ap_return_8;
output  [31:0] ap_return_9;
output  [31:0] ap_return_10;
output  [31:0] ap_return_11;
output  [31:0] ap_return_12;
output  [31:0] ap_return_13;
output  [31:0] ap_return_14;
output  [31:0] ap_return_15;
output  [31:0] ap_return_16;
output  [31:0] ap_return_17;
output  [31:0] ap_return_18;
output  [31:0] ap_return_19;
output  [31:0] ap_return_20;
output  [31:0] ap_return_21;
output  [31:0] ap_return_22;
output  [31:0] ap_return_23;
output  [31:0] ap_return_24;
output  [31:0] ap_return_25;
output  [31:0] ap_return_26;
output  [31:0] ap_return_27;
output  [31:0] ap_return_28;
output  [31:0] ap_return_29;
output  [31:0] ap_return_30;
output  [31:0] ap_return_31;
wire tmp_0_3;
assign tmp_0_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]);
wire tmp_0_7;
assign tmp_0_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]);
wire tmp_0_8;
assign tmp_0_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]);
wire tmp_0_11;
assign tmp_0_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]);
wire tmp_0_13;
assign tmp_0_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]);
wire tmp_0_14;
assign tmp_0_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]);
wire tmp_0_16;
assign tmp_0_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]);
wire tmp_0_18;
assign tmp_0_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]);
wire tmp_0_19;
assign tmp_0_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]);
wire tmp_0_21;
assign tmp_0_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]);
wire tmp_0_25;
assign tmp_0_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]);
wire tmp_0_27;
assign tmp_0_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]);
wire tmp_0_28;
assign tmp_0_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]);
wire tmp_0_31;
assign tmp_0_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]);
assign ap_return_0 = {1'b0,1'b0,1'b0,tmp_0_3,1'b0,1'b0,1'b0,tmp_0_7,tmp_0_8,1'b0,1'b0,tmp_0_11,1'b0,tmp_0_13,tmp_0_14,1'b0,tmp_0_16,1'b0,tmp_0_18,tmp_0_19,1'b0,tmp_0_21,1'b0,1'b0,1'b0,tmp_0_25,1'b0,tmp_0_27,tmp_0_28,1'b0,1'b0,tmp_0_31};
wire tmp_1_0;
assign tmp_1_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]);
wire tmp_1_7;
assign tmp_1_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]);
wire tmp_1_10;
assign tmp_1_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]);
wire tmp_1_13;
assign tmp_1_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]);
wire tmp_1_15;
assign tmp_1_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]);
wire tmp_1_16;
assign tmp_1_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]);
wire tmp_1_18;
assign tmp_1_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]);
wire tmp_1_21;
assign tmp_1_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]);
wire tmp_1_29;
assign tmp_1_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]);
wire tmp_1_30;
assign tmp_1_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]);
wire tmp_1_31;
assign tmp_1_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]);
assign ap_return_1 = {tmp_1_0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_1_7,1'b0,1'b0,tmp_1_10,1'b0,1'b0,tmp_1_13,1'b0,tmp_1_15,tmp_1_16,1'b0,tmp_1_18,1'b0,1'b0,tmp_1_21,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_1_29,tmp_1_30,tmp_1_31};
wire tmp_2_3;
assign tmp_2_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]);
wire tmp_2_16;
assign tmp_2_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]);
wire tmp_2_23;
assign tmp_2_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]);
wire tmp_2_31;
assign tmp_2_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]);
assign ap_return_2 = {1'b0,1'b0,1'b0,tmp_2_3,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_2_16,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_2_23,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_2_31};
wire tmp_3_3;
assign tmp_3_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]);
wire tmp_3_16;
assign tmp_3_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]);
wire tmp_3_17;
assign tmp_3_17 = (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]);
wire tmp_3_22;
assign tmp_3_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]);
wire tmp_3_26;
assign tmp_3_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]);
wire tmp_3_29;
assign tmp_3_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]);
wire tmp_3_30;
assign tmp_3_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]);
wire tmp_3_31;
assign tmp_3_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]);
assign ap_return_3 = {1'b0,1'b0,1'b0,tmp_3_3,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_3_16,tmp_3_17,1'b0,1'b0,1'b0,1'b0,tmp_3_22,1'b0,1'b0,1'b0,tmp_3_26,1'b0,1'b0,tmp_3_29,tmp_3_30,tmp_3_31};
wire tmp_4_0;
assign tmp_4_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]);
wire tmp_4_14;
assign tmp_4_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]);
wire tmp_4_16;
assign tmp_4_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]);
wire tmp_4_18;
assign tmp_4_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]);
wire tmp_4_21;
assign tmp_4_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]);
wire tmp_4_29;
assign tmp_4_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]);
assign ap_return_4 = {tmp_4_0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_4_14,1'b0,tmp_4_16,1'b0,tmp_4_18,1'b0,1'b0,tmp_4_21,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_4_29,1'b0,1'b0};
wire tmp_5_0;
assign tmp_5_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]);
wire tmp_5_3;
assign tmp_5_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]);
wire tmp_5_4;
assign tmp_5_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]);
wire tmp_5_7;
assign tmp_5_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]);
wire tmp_5_10;
assign tmp_5_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]);
wire tmp_5_13;
assign tmp_5_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]);
wire tmp_5_14;
assign tmp_5_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]);
wire tmp_5_16;
assign tmp_5_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]);
wire tmp_5_17;
assign tmp_5_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]);
wire tmp_5_18;
assign tmp_5_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]);
wire tmp_5_21;
assign tmp_5_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]);
wire tmp_5_24;
assign tmp_5_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]);
wire tmp_5_29;
assign tmp_5_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]);
wire tmp_5_30;
assign tmp_5_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]);
wire tmp_5_31;
assign tmp_5_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]);
assign ap_return_5 = {tmp_5_0,1'b0,1'b0,tmp_5_3,tmp_5_4,1'b0,1'b0,tmp_5_7,1'b0,1'b0,tmp_5_10,1'b0,1'b0,tmp_5_13,tmp_5_14,1'b0,tmp_5_16,tmp_5_17,tmp_5_18,1'b0,1'b0,tmp_5_21,1'b0,1'b0,tmp_5_24,1'b0,1'b0,1'b0,1'b0,tmp_5_29,tmp_5_30,tmp_5_31};
wire tmp_6_3;
assign tmp_6_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]);
wire tmp_6_5;
assign tmp_6_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]);
wire tmp_6_7;
assign tmp_6_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]);
wire tmp_6_9;
assign tmp_6_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]);
wire tmp_6_16;
assign tmp_6_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]);
wire tmp_6_17;
assign tmp_6_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]);
wire tmp_6_22;
assign tmp_6_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]);
wire tmp_6_23;
assign tmp_6_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]);
wire tmp_6_29;
assign tmp_6_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]);
wire tmp_6_30;
assign tmp_6_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]);
wire tmp_6_31;
assign tmp_6_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]);
assign ap_return_6 = {1'b0,1'b0,1'b0,tmp_6_3,1'b0,tmp_6_5,1'b0,tmp_6_7,1'b0,tmp_6_9,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_6_16,tmp_6_17,1'b0,1'b0,1'b0,1'b0,tmp_6_22,tmp_6_23,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_6_29,tmp_6_30,tmp_6_31};
wire tmp_7_3;
assign tmp_7_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]);
wire tmp_7_7;
assign tmp_7_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]);
wire tmp_7_16;
assign tmp_7_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]);
wire tmp_7_21;
assign tmp_7_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]);
wire tmp_7_26;
assign tmp_7_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]);
wire tmp_7_29;
assign tmp_7_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]);
wire tmp_7_31;
assign tmp_7_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]);
assign ap_return_7 = {1'b0,1'b0,1'b0,tmp_7_3,1'b0,1'b0,1'b0,tmp_7_7,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_7_16,1'b0,1'b0,1'b0,1'b0,tmp_7_21,1'b0,1'b0,1'b0,1'b0,tmp_7_26,1'b0,1'b0,tmp_7_29,1'b0,tmp_7_31};
wire tmp_8_0;
assign tmp_8_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]);
wire tmp_8_3;
assign tmp_8_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]);
wire tmp_8_6;
assign tmp_8_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]);
wire tmp_8_17;
assign tmp_8_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]);
wire tmp_8_23;
assign tmp_8_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]);
wire tmp_8_24;
assign tmp_8_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]);
wire tmp_8_29;
assign tmp_8_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]);
wire tmp_8_31;
assign tmp_8_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_8_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_8_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_8_V_read[31]);
assign ap_return_8 = {tmp_8_0,1'b0,1'b0,tmp_8_3,1'b0,1'b0,tmp_8_6,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_8_17,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_8_23,tmp_8_24,1'b0,1'b0,1'b0,1'b0,tmp_8_29,1'b0,tmp_8_31};
wire tmp_9_0;
assign tmp_9_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]);
wire tmp_9_3;
assign tmp_9_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]);
wire tmp_9_16;
assign tmp_9_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]);
wire tmp_9_17;
assign tmp_9_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]);
wire tmp_9_18;
assign tmp_9_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]);
wire tmp_9_20;
assign tmp_9_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]);
wire tmp_9_21;
assign tmp_9_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]);
wire tmp_9_22;
assign tmp_9_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]);
wire tmp_9_23;
assign tmp_9_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]);
wire tmp_9_24;
assign tmp_9_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]);
wire tmp_9_31;
assign tmp_9_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]);
assign ap_return_9 = {tmp_9_0,1'b0,1'b0,tmp_9_3,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_9_16,tmp_9_17,tmp_9_18,1'b0,tmp_9_20,tmp_9_21,tmp_9_22,tmp_9_23,tmp_9_24,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_9_31};
wire tmp_10_21;
assign tmp_10_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]);
wire tmp_10_26;
assign tmp_10_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]);
wire tmp_10_29;
assign tmp_10_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]);
wire tmp_10_31;
assign tmp_10_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]);
assign ap_return_10 = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_10_21,1'b0,1'b0,1'b0,1'b0,tmp_10_26,1'b0,1'b0,tmp_10_29,1'b0,tmp_10_31};
wire tmp_11_3;
assign tmp_11_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]);
wire tmp_11_17;
assign tmp_11_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]);
wire tmp_11_20;
assign tmp_11_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]);
wire tmp_11_21;
assign tmp_11_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]);
wire tmp_11_24;
assign tmp_11_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]);
wire tmp_11_26;
assign tmp_11_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]);
wire tmp_11_29;
assign tmp_11_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]);
wire tmp_11_30;
assign tmp_11_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]);
assign ap_return_11 = {1'b0,1'b0,1'b0,tmp_11_3,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_11_17,1'b0,1'b0,tmp_11_20,tmp_11_21,1'b0,1'b0,tmp_11_24,1'b0,tmp_11_26,1'b0,1'b0,tmp_11_29,tmp_11_30,1'b0};
wire tmp_12_0;
assign tmp_12_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]);
wire tmp_12_3;
assign tmp_12_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]);
wire tmp_12_6;
assign tmp_12_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]);
wire tmp_12_9;
assign tmp_12_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]);
wire tmp_12_13;
assign tmp_12_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]);
wire tmp_12_17;
assign tmp_12_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]);
wire tmp_12_19;
assign tmp_12_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]);
wire tmp_12_23;
assign tmp_12_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]);
wire tmp_12_24;
assign tmp_12_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]);
wire tmp_12_25;
assign tmp_12_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]);
wire tmp_12_29;
assign tmp_12_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]);
wire tmp_12_31;
assign tmp_12_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]);
assign ap_return_12 = {tmp_12_0,1'b0,1'b0,tmp_12_3,1'b0,1'b0,tmp_12_6,1'b0,1'b0,tmp_12_9,1'b0,1'b0,1'b0,tmp_12_13,1'b0,1'b0,1'b0,tmp_12_17,1'b0,tmp_12_19,1'b0,1'b0,1'b0,tmp_12_23,tmp_12_24,tmp_12_25,1'b0,1'b0,1'b0,tmp_12_29,1'b0,tmp_12_31};
wire tmp_13_3;
assign tmp_13_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]);
wire tmp_13_7;
assign tmp_13_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]);
wire tmp_13_8;
assign tmp_13_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]);
wire tmp_13_13;
assign tmp_13_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]);
wire tmp_13_16;
assign tmp_13_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]);
wire tmp_13_19;
assign tmp_13_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]);
wire tmp_13_21;
assign tmp_13_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]);
wire tmp_13_22;
assign tmp_13_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]);
wire tmp_13_27;
assign tmp_13_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]);
wire tmp_13_30;
assign tmp_13_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]);
wire tmp_13_31;
assign tmp_13_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]);
assign ap_return_13 = {1'b0,1'b0,1'b0,tmp_13_3,1'b0,1'b0,1'b0,tmp_13_7,tmp_13_8,1'b0,1'b0,1'b0,1'b0,tmp_13_13,1'b0,1'b0,tmp_13_16,1'b0,1'b0,tmp_13_19,1'b0,tmp_13_21,tmp_13_22,1'b0,1'b0,1'b0,1'b0,tmp_13_27,1'b0,1'b0,tmp_13_30,tmp_13_31};
wire tmp_14_0;
assign tmp_14_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]);
wire tmp_14_16;
assign tmp_14_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]);
wire tmp_14_17;
assign tmp_14_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]);
wire tmp_14_18;
assign tmp_14_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]);
wire tmp_14_21;
assign tmp_14_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]);
wire tmp_14_23;
assign tmp_14_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]);
assign ap_return_14 = {tmp_14_0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_14_16,tmp_14_17,tmp_14_18,1'b0,1'b0,tmp_14_21,1'b0,tmp_14_23,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
wire tmp_15_3;
assign tmp_15_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]);
wire tmp_15_7;
assign tmp_15_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]);
wire tmp_15_9;
assign tmp_15_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]);
wire tmp_15_18;
assign tmp_15_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]);
wire tmp_15_19;
assign tmp_15_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]);
wire tmp_15_20;
assign tmp_15_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]);
wire tmp_15_21;
assign tmp_15_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]);
wire tmp_15_23;
assign tmp_15_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]);
wire tmp_15_24;
assign tmp_15_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]);
wire tmp_15_29;
assign tmp_15_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]);
wire tmp_15_31;
assign tmp_15_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_15_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_15_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_15_V_read[31]);
assign ap_return_15 = {1'b0,1'b0,1'b0,tmp_15_3,1'b0,1'b0,1'b0,tmp_15_7,1'b0,tmp_15_9,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_15_18,tmp_15_19,tmp_15_20,tmp_15_21,1'b0,tmp_15_23,tmp_15_24,1'b0,1'b0,1'b0,1'b0,tmp_15_29,1'b0,tmp_15_31};
wire tmp_16_0;
assign tmp_16_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_16_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_16_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_16_V_read[0]);
wire tmp_16_3;
assign tmp_16_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_16_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_16_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_16_V_read[3]);
wire tmp_16_11;
assign tmp_16_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_16_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_16_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_16_V_read[11]);
wire tmp_16_18;
assign tmp_16_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_16_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_16_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_16_V_read[18]);
wire tmp_16_19;
assign tmp_16_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_16_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_16_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_16_V_read[19]);
wire tmp_16_21;
assign tmp_16_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_16_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_16_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_16_V_read[21]);
wire tmp_16_23;
assign tmp_16_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_16_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_16_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_16_V_read[23]);
wire tmp_16_24;
assign tmp_16_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_16_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_16_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_16_V_read[24]);
wire tmp_16_29;
assign tmp_16_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_16_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_16_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_16_V_read[29]);
wire tmp_16_31;
assign tmp_16_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_16_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_16_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_16_V_read[31]);
assign ap_return_16 = {tmp_16_0,1'b0,1'b0,tmp_16_3,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_16_11,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_16_18,tmp_16_19,1'b0,tmp_16_21,1'b0,tmp_16_23,tmp_16_24,1'b0,1'b0,1'b0,1'b0,tmp_16_29,1'b0,tmp_16_31};
wire tmp_17_0;
assign tmp_17_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_17_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_17_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_17_V_read[0]);
wire tmp_17_3;
assign tmp_17_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_17_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_17_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_17_V_read[3]);
wire tmp_17_5;
assign tmp_17_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_17_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_17_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_17_V_read[5]);
wire tmp_17_8;
assign tmp_17_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_17_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_17_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_17_V_read[8]);
wire tmp_17_17;
assign tmp_17_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_17_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_17_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_17_V_read[17]);
wire tmp_17_19;
assign tmp_17_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_17_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_17_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_17_V_read[19]);
wire tmp_17_21;
assign tmp_17_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_17_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_17_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_17_V_read[21]);
wire tmp_17_22;
assign tmp_17_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_17_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_17_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_17_V_read[22]);
assign ap_return_17 = {tmp_17_0,1'b0,1'b0,tmp_17_3,1'b0,tmp_17_5,1'b0,1'b0,tmp_17_8,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_17_17,1'b0,tmp_17_19,1'b0,tmp_17_21,tmp_17_22,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
wire tmp_18_0;
assign tmp_18_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_18_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_18_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_18_V_read[0]);
wire tmp_18_7;
assign tmp_18_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_18_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_18_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_18_V_read[7]);
wire tmp_18_10;
assign tmp_18_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_18_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_18_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_18_V_read[10]);
wire tmp_18_16;
assign tmp_18_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_18_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_18_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_18_V_read[16]);
wire tmp_18_17;
assign tmp_18_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_18_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_18_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_18_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_18_V_read[17]);
wire tmp_18_19;
assign tmp_18_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_18_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_18_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_18_V_read[19]);
wire tmp_18_23;
assign tmp_18_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_18_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_18_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_18_V_read[23]);
wire tmp_18_25;
assign tmp_18_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_18_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_18_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_18_V_read[25]);
wire tmp_18_29;
assign tmp_18_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_18_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_18_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_18_V_read[29]);
wire tmp_18_31;
assign tmp_18_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_18_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_18_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_18_V_read[31]);
assign ap_return_18 = {tmp_18_0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_18_7,1'b0,1'b0,tmp_18_10,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_18_16,tmp_18_17,1'b0,tmp_18_19,1'b0,1'b0,1'b0,tmp_18_23,1'b0,tmp_18_25,1'b0,1'b0,1'b0,tmp_18_29,1'b0,tmp_18_31};
wire tmp_19_7;
assign tmp_19_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_19_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_19_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_19_V_read[7]);
wire tmp_19_12;
assign tmp_19_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_19_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_19_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_19_V_read[12]);
wire tmp_19_16;
assign tmp_19_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_19_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_19_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_19_V_read[16]);
wire tmp_19_22;
assign tmp_19_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_19_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_19_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_19_V_read[22]);
wire tmp_19_26;
assign tmp_19_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_19_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_19_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_19_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_19_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_19_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_19_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_19_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_19_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_19_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_19_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_19_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_19_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_19_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_19_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_19_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_19_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_19_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_19_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_19_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_19_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_19_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_19_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_19_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_19_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_19_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_19_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_19_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_19_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_19_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_19_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_19_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_19_V_read[26]);
assign ap_return_19 = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_19_7,1'b0,1'b0,1'b0,1'b0,tmp_19_12,1'b0,1'b0,1'b0,tmp_19_16,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_19_22,1'b0,1'b0,1'b0,tmp_19_26,1'b0,1'b0,1'b0,1'b0,1'b0};
wire tmp_20_0;
assign tmp_20_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_20_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_20_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_20_V_read[0]);
wire tmp_20_3;
assign tmp_20_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_20_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_20_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_20_V_read[3]);
wire tmp_20_5;
assign tmp_20_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_20_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_20_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_20_V_read[5]);
wire tmp_20_8;
assign tmp_20_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_20_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_20_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_20_V_read[8]);
wire tmp_20_16;
assign tmp_20_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_20_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_20_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_20_V_read[16]);
wire tmp_20_17;
assign tmp_20_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_20_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_20_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_20_V_read[17]);
wire tmp_20_21;
assign tmp_20_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_20_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_20_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_20_V_read[21]);
wire tmp_20_28;
assign tmp_20_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_20_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_20_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_20_V_read[28]);
assign ap_return_20 = {tmp_20_0,1'b0,1'b0,tmp_20_3,1'b0,tmp_20_5,1'b0,1'b0,tmp_20_8,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_20_16,tmp_20_17,1'b0,1'b0,1'b0,tmp_20_21,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_20_28,1'b0,1'b0,1'b0};
wire tmp_21_0;
assign tmp_21_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_21_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_21_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_21_V_read[0]);
wire tmp_21_7;
assign tmp_21_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_21_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_21_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_21_V_read[7]);
wire tmp_21_8;
assign tmp_21_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_21_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_21_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_21_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_21_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_21_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_21_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_21_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_21_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_21_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_21_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_21_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_21_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_21_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_21_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_21_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_21_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_21_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_21_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_21_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_21_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_21_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_21_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_21_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_21_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_21_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_21_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_21_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_21_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_21_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_21_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_21_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_21_V_read[8]);
wire tmp_21_16;
assign tmp_21_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_21_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_21_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_21_V_read[16]);
wire tmp_21_21;
assign tmp_21_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_21_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_21_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_21_V_read[21]);
wire tmp_21_24;
assign tmp_21_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_21_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_21_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_21_V_read[24]);
wire tmp_21_26;
assign tmp_21_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_21_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_21_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_21_V_read[26]);
wire tmp_21_28;
assign tmp_21_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_21_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_21_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_21_V_read[28]);
wire tmp_21_29;
assign tmp_21_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_21_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_21_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_21_V_read[29]);
wire tmp_21_30;
assign tmp_21_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_21_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_21_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_21_V_read[30]);
wire tmp_21_31;
assign tmp_21_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_21_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_21_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_21_V_read[31]);
assign ap_return_21 = {tmp_21_0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_21_7,tmp_21_8,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_21_16,1'b0,1'b0,1'b0,1'b0,tmp_21_21,1'b0,1'b0,tmp_21_24,1'b0,tmp_21_26,1'b0,tmp_21_28,tmp_21_29,tmp_21_30,tmp_21_31};
wire tmp_22_0;
assign tmp_22_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_22_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_22_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_22_V_read[0]);
wire tmp_22_1;
assign tmp_22_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_22_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_22_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_22_V_read[1]);
wire tmp_22_3;
assign tmp_22_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_22_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_22_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_22_V_read[3]);
wire tmp_22_6;
assign tmp_22_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_22_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_22_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_22_V_read[6]);
wire tmp_22_8;
assign tmp_22_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_22_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_22_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_22_V_read[8]);
wire tmp_22_17;
assign tmp_22_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_22_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_22_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_22_V_read[17]);
wire tmp_22_21;
assign tmp_22_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_22_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_22_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_22_V_read[21]);
wire tmp_22_22;
assign tmp_22_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_22_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_22_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_22_V_read[22]);
wire tmp_22_23;
assign tmp_22_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_22_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_22_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_22_V_read[23]);
wire tmp_22_26;
assign tmp_22_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_22_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_22_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_22_V_read[26]);
wire tmp_22_29;
assign tmp_22_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_22_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_22_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_22_V_read[29]);
wire tmp_22_31;
assign tmp_22_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_22_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_22_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_22_V_read[31]);
assign ap_return_22 = {tmp_22_0,tmp_22_1,1'b0,tmp_22_3,1'b0,1'b0,tmp_22_6,1'b0,tmp_22_8,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_22_17,1'b0,1'b0,1'b0,tmp_22_21,tmp_22_22,tmp_22_23,1'b0,1'b0,tmp_22_26,1'b0,1'b0,tmp_22_29,1'b0,tmp_22_31};
wire tmp_23_0;
assign tmp_23_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_23_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_23_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_23_V_read[0]);
wire tmp_23_1;
assign tmp_23_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_23_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_23_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_23_V_read[1]);
wire tmp_23_7;
assign tmp_23_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_23_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_23_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_23_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_23_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_23_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_23_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_23_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_23_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_23_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_23_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_23_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_23_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_23_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_23_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_23_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_23_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_23_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_23_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_23_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_23_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_23_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_23_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_23_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_23_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_23_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_23_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_23_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_23_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_23_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_23_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_23_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_23_V_read[7]);
wire tmp_23_15;
assign tmp_23_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_23_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_23_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_23_V_read[15]);
wire tmp_23_17;
assign tmp_23_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_23_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_23_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_23_V_read[17]);
wire tmp_23_18;
assign tmp_23_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_23_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_23_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_23_V_read[18]);
wire tmp_23_26;
assign tmp_23_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_23_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_23_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_23_V_read[26]);
wire tmp_23_29;
assign tmp_23_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_23_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_23_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_23_V_read[29]);
assign ap_return_23 = {tmp_23_0,tmp_23_1,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_23_7,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_23_15,1'b0,tmp_23_17,tmp_23_18,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_23_26,1'b0,1'b0,tmp_23_29,1'b0,1'b0};
wire tmp_24_0;
assign tmp_24_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_24_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_24_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_24_V_read[0]);
wire tmp_24_8;
assign tmp_24_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_24_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_24_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_24_V_read[8]);
wire tmp_24_16;
assign tmp_24_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_24_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_24_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_24_V_read[16]);
wire tmp_24_23;
assign tmp_24_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_24_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_24_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_24_V_read[23]);
wire tmp_24_27;
assign tmp_24_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_24_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_24_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_24_V_read[27]);
wire tmp_24_29;
assign tmp_24_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_24_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_24_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_24_V_read[29]);
wire tmp_24_31;
assign tmp_24_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_24_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_24_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_24_V_read[31]);
assign ap_return_24 = {tmp_24_0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_24_8,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_24_16,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_24_23,1'b0,1'b0,1'b0,tmp_24_27,1'b0,tmp_24_29,1'b0,tmp_24_31};
wire tmp_25_8;
assign tmp_25_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_25_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_25_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_25_V_read[8]);
wire tmp_25_13;
assign tmp_25_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_25_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_25_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_25_V_read[13]);
wire tmp_25_21;
assign tmp_25_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_25_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_25_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_25_V_read[21]);
wire tmp_25_24;
assign tmp_25_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_25_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_25_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_25_V_read[24]);
wire tmp_25_29;
assign tmp_25_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_25_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_25_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_25_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_25_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_25_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_25_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_25_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_25_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_25_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_25_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_25_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_25_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_25_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_25_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_25_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_25_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_25_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_25_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_25_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_25_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_25_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_25_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_25_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_25_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_25_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_25_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_25_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_25_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_25_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_25_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_25_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_25_V_read[29]);
assign ap_return_25 = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_25_8,1'b0,1'b0,1'b0,1'b0,tmp_25_13,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_25_21,1'b0,1'b0,tmp_25_24,1'b0,1'b0,1'b0,1'b0,tmp_25_29,1'b0,1'b0};
wire tmp_26_2;
assign tmp_26_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_26_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_26_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_26_V_read[2]);
wire tmp_26_9;
assign tmp_26_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_26_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_26_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_26_V_read[9]);
wire tmp_26_16;
assign tmp_26_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_26_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_26_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_26_V_read[16]);
wire tmp_26_17;
assign tmp_26_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_26_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_26_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_26_V_read[17]);
wire tmp_26_23;
assign tmp_26_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_26_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_26_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_26_V_read[23]);
wire tmp_26_24;
assign tmp_26_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_26_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_26_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_26_V_read[24]);
wire tmp_26_29;
assign tmp_26_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_26_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_26_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_26_V_read[29]);
assign ap_return_26 = {1'b0,1'b0,tmp_26_2,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_26_9,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_26_16,tmp_26_17,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_26_23,tmp_26_24,1'b0,1'b0,1'b0,1'b0,tmp_26_29,1'b0,1'b0};
wire tmp_27_2;
assign tmp_27_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_27_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_27_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_27_V_read[2]);
wire tmp_27_5;
assign tmp_27_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_27_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_27_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_27_V_read[5]);
wire tmp_27_7;
assign tmp_27_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_27_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_27_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_27_V_read[7]);
wire tmp_27_14;
assign tmp_27_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_27_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_27_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_27_V_read[14]);
wire tmp_27_16;
assign tmp_27_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_27_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_27_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_27_V_read[16]);
wire tmp_27_21;
assign tmp_27_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_27_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_27_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_27_V_read[21]);
wire tmp_27_25;
assign tmp_27_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_27_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_27_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_27_V_read[25]);
wire tmp_27_31;
assign tmp_27_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_27_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_27_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_27_V_read[31]);
assign ap_return_27 = {1'b0,1'b0,tmp_27_2,1'b0,1'b0,tmp_27_5,1'b0,tmp_27_7,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_27_14,1'b0,tmp_27_16,1'b0,1'b0,1'b0,1'b0,tmp_27_21,1'b0,1'b0,1'b0,tmp_27_25,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_27_31};
wire tmp_28_0;
assign tmp_28_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_28_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_28_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_28_V_read[0]);
wire tmp_28_3;
assign tmp_28_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_28_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_28_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_28_V_read[3]);
wire tmp_28_7;
assign tmp_28_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_28_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_28_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_28_V_read[7]);
wire tmp_28_13;
assign tmp_28_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_28_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_28_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_28_V_read[13]);
wire tmp_28_16;
assign tmp_28_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_28_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_28_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_28_V_read[16]);
wire tmp_28_21;
assign tmp_28_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_28_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_28_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_28_V_read[21]);
wire tmp_28_24;
assign tmp_28_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_28_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_28_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_28_V_read[24]);
wire tmp_28_26;
assign tmp_28_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_28_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_28_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_28_V_read[26]);
wire tmp_28_28;
assign tmp_28_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_28_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_28_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_28_V_read[28]);
wire tmp_28_30;
assign tmp_28_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_28_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_28_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_28_V_read[30]);
wire tmp_28_31;
assign tmp_28_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_28_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_28_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_28_V_read[31]);
assign ap_return_28 = {tmp_28_0,1'b0,1'b0,tmp_28_3,1'b0,1'b0,1'b0,tmp_28_7,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_28_13,1'b0,1'b0,tmp_28_16,1'b0,1'b0,1'b0,1'b0,tmp_28_21,1'b0,1'b0,tmp_28_24,1'b0,tmp_28_26,1'b0,tmp_28_28,1'b0,tmp_28_30,tmp_28_31};
wire tmp_29_0;
assign tmp_29_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_29_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_29_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_29_V_read[0]);
wire tmp_29_7;
assign tmp_29_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_29_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_29_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_29_V_read[7]);
wire tmp_29_11;
assign tmp_29_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_29_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_29_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_29_V_read[11]);
wire tmp_29_16;
assign tmp_29_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_29_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_29_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_29_V_read[16]);
wire tmp_29_17;
assign tmp_29_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_29_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_29_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_29_V_read[17]);
wire tmp_29_22;
assign tmp_29_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_29_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_29_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_29_V_read[22]);
wire tmp_29_23;
assign tmp_29_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_29_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_29_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_29_V_read[23]);
wire tmp_29_25;
assign tmp_29_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_29_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_29_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_29_V_read[25]);
wire tmp_29_29;
assign tmp_29_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_29_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_29_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_29_V_read[29]);
wire tmp_29_30;
assign tmp_29_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_29_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_29_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_29_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_29_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_29_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_29_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_29_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_29_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_29_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_29_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_29_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_29_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_29_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_29_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_29_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_29_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_29_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_29_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_29_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_29_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_29_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_29_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_29_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_29_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_29_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_29_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_29_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_29_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_29_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_29_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_29_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_29_V_read[30]);
assign ap_return_29 = {tmp_29_0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_29_7,1'b0,1'b0,1'b0,tmp_29_11,1'b0,1'b0,1'b0,1'b0,tmp_29_16,tmp_29_17,1'b0,1'b0,1'b0,1'b0,tmp_29_22,tmp_29_23,1'b0,tmp_29_25,1'b0,1'b0,1'b0,tmp_29_29,tmp_29_30,1'b0};
wire tmp_30_0;
assign tmp_30_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_30_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_30_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_30_V_read[0]);
wire tmp_30_3;
assign tmp_30_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_30_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_30_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_30_V_read[3]);
wire tmp_30_6;
assign tmp_30_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_30_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_30_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_30_V_read[6]);
wire tmp_30_8;
assign tmp_30_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_30_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_30_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_30_V_read[8]);
wire tmp_30_9;
assign tmp_30_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_30_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_30_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_30_V_read[9]);
wire tmp_30_10;
assign tmp_30_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_30_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_30_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_30_V_read[10]);
wire tmp_30_11;
assign tmp_30_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_30_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_30_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_30_V_read[11]);
wire tmp_30_19;
assign tmp_30_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_30_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_30_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_30_V_read[19]);
wire tmp_30_21;
assign tmp_30_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_30_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_30_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_30_V_read[21]);
wire tmp_30_24;
assign tmp_30_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_30_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_30_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_30_V_read[24]);
wire tmp_30_25;
assign tmp_30_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_30_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_30_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_30_V_read[25]);
wire tmp_30_31;
assign tmp_30_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_30_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_30_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_30_V_read[31]);
assign ap_return_30 = {tmp_30_0,1'b0,1'b0,tmp_30_3,1'b0,1'b0,tmp_30_6,1'b0,tmp_30_8,tmp_30_9,tmp_30_10,tmp_30_11,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_30_19,1'b0,tmp_30_21,1'b0,1'b0,tmp_30_24,tmp_30_25,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_30_31};
wire tmp_31_0;
assign tmp_31_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_31_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_31_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_31_V_read[0]);
wire tmp_31_3;
assign tmp_31_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_31_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_31_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_31_V_read[3]);
wire tmp_31_7;
assign tmp_31_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_31_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_31_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_31_V_read[7]);
wire tmp_31_8;
assign tmp_31_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_31_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_31_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_31_V_read[8]);
wire tmp_31_23;
assign tmp_31_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_31_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_31_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_31_V_read[23]);
wire tmp_31_28;
assign tmp_31_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_31_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_31_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_31_V_read[28]);
wire tmp_31_29;
assign tmp_31_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_31_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_31_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_31_V_read[29]);
wire tmp_31_31;
assign tmp_31_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_31_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_31_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_31_V_read[31]);
assign ap_return_31 = {tmp_31_0,1'b0,1'b0,tmp_31_3,1'b0,1'b0,1'b0,tmp_31_7,tmp_31_8,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,tmp_31_23,1'b0,1'b0,1'b0,1'b0,tmp_31_28,tmp_31_29,1'b0,tmp_31_31};
endmodule