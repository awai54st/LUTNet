`timescale 1 ns / 1 ps

module LUTARRAY_36u_4u_s (
        in_V,
        in_1_V,
        in_2_V,
        in_3_V,
        weight_0_0_V_read,
        weight_0_1_V_read,
        weight_0_2_V_read,
        weight_0_3_V_read,
        weight_0_4_V_read,
        weight_0_5_V_read,
        weight_0_6_V_read,
        weight_0_7_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7);



input  [71:0] in_V;
input  [71:0] in_1_V;
input  [71:0] in_2_V;
input  [71:0] in_3_V;
input  [95:0] weight_0_0_V_read;
input  [95:0] weight_0_1_V_read;
input  [95:0] weight_0_2_V_read;
input  [95:0] weight_0_3_V_read;
input  [95:0] weight_0_4_V_read;
input  [95:0] weight_0_5_V_read;
input  [95:0] weight_0_6_V_read;
input  [95:0] weight_0_7_V_read;
output  [71:0] ap_return_0;
output  [71:0] ap_return_1;
output  [71:0] ap_return_2;
output  [71:0] ap_return_3;
output  [71:0] ap_return_4;
output  [71:0] ap_return_5;
output  [71:0] ap_return_6;
output  [71:0] ap_return_7;
wire tmp_0_0;
assign tmp_0_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_0_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_0_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_0_V_read[0]);
wire tmp_0_1;
assign tmp_0_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]);
wire tmp_0_2;
assign tmp_0_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]);
wire tmp_0_3;
assign tmp_0_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]);
wire tmp_0_4;
assign tmp_0_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]);
wire tmp_0_6;
assign tmp_0_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]);
wire tmp_0_7;
assign tmp_0_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_0_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_0_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_0_V_read[7]);
wire tmp_0_8;
assign tmp_0_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]);
wire tmp_0_9;
assign tmp_0_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_0_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_0_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_0_V_read[9]);
wire tmp_0_10;
assign tmp_0_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]);
wire tmp_0_11;
assign tmp_0_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]);
wire tmp_0_12;
assign tmp_0_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]);
wire tmp_0_13;
assign tmp_0_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]);
wire tmp_0_14;
assign tmp_0_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]);
wire tmp_0_15;
assign tmp_0_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]);
wire tmp_0_16;
assign tmp_0_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]);
wire tmp_0_17;
assign tmp_0_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]);
wire tmp_0_18;
assign tmp_0_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]);
wire tmp_0_19;
assign tmp_0_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]);
wire tmp_0_20;
assign tmp_0_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]);
wire tmp_0_21;
assign tmp_0_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]);
wire tmp_0_22;
assign tmp_0_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]);
wire tmp_0_23;
assign tmp_0_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]);
wire tmp_0_24;
assign tmp_0_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]);
wire tmp_0_25;
assign tmp_0_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]);
wire tmp_0_26;
assign tmp_0_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_0_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_0_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_0_V_read[26]);
wire tmp_0_27;
assign tmp_0_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]);
wire tmp_0_28;
assign tmp_0_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]);
wire tmp_0_29;
assign tmp_0_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_0_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_0_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_0_V_read[29]);
wire tmp_0_30;
assign tmp_0_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]);
wire tmp_0_31;
assign tmp_0_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_0_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_0_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_0_V_read[31]);
wire tmp_0_32;
assign tmp_0_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]);
wire tmp_0_33;
assign tmp_0_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]);
wire tmp_0_34;
assign tmp_0_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]);
wire tmp_0_35;
assign tmp_0_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]);
wire tmp_0_36;
assign tmp_0_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]);
wire tmp_0_37;
assign tmp_0_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]);
wire tmp_0_38;
assign tmp_0_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_0_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_0_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_0_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_0_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_0_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_0_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_0_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_0_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_0_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_0_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_0_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_0_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_0_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_0_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_0_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_0_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_0_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_0_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_0_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_0_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_0_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_0_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_0_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_0_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_0_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_0_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_0_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_0_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_0_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_0_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_0_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_0_V_read[38]);
wire tmp_0_39;
assign tmp_0_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_0_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_0_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_0_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_0_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_0_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_0_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_0_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_0_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_0_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_0_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_0_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_0_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_0_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_0_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_0_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_0_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_0_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_0_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_0_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_0_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_0_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_0_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_0_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_0_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_0_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_0_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_0_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_0_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_0_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_0_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_0_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_0_V_read[39]);
wire tmp_0_40;
assign tmp_0_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]);
wire tmp_0_41;
assign tmp_0_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]);
wire tmp_0_42;
assign tmp_0_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]);
wire tmp_0_43;
assign tmp_0_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]);
wire tmp_0_44;
assign tmp_0_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]);
wire tmp_0_45;
assign tmp_0_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]);
wire tmp_0_46;
assign tmp_0_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]);
wire tmp_0_47;
assign tmp_0_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_0_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_0_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_0_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_0_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_0_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_0_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_0_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_0_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_0_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_0_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_0_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_0_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_0_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_0_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_0_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_0_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_0_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_0_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_0_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_0_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_0_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_0_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_0_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_0_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_0_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_0_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_0_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_0_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_0_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_0_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_0_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_0_V_read[47]);
wire tmp_0_48;
assign tmp_0_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]);
wire tmp_0_49;
assign tmp_0_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]);
wire tmp_0_50;
assign tmp_0_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]);
wire tmp_0_51;
assign tmp_0_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]);
wire tmp_0_52;
assign tmp_0_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]);
wire tmp_0_53;
assign tmp_0_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]);
wire tmp_0_54;
assign tmp_0_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]);
wire tmp_0_55;
assign tmp_0_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]);
wire tmp_0_56;
assign tmp_0_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]);
wire tmp_0_57;
assign tmp_0_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]);
wire tmp_0_58;
assign tmp_0_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]);
wire tmp_0_59;
assign tmp_0_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]);
wire tmp_0_60;
assign tmp_0_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]);
wire tmp_0_61;
assign tmp_0_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]);
wire tmp_0_62;
assign tmp_0_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]);
wire tmp_0_63;
assign tmp_0_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]);
wire tmp_0_64;
assign tmp_0_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]);
wire tmp_0_65;
assign tmp_0_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]);
wire tmp_0_66;
assign tmp_0_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]);
wire tmp_0_67;
assign tmp_0_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]);
wire tmp_0_68;
assign tmp_0_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]);
wire tmp_0_69;
assign tmp_0_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]);
wire tmp_0_70;
assign tmp_0_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]);
wire tmp_0_71;
assign tmp_0_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]);
assign ap_return_0 = {tmp_0_0,tmp_0_1,tmp_0_2,tmp_0_3,tmp_0_4,1'b0,tmp_0_6,tmp_0_7,tmp_0_8,tmp_0_9,tmp_0_10,tmp_0_11,tmp_0_12,tmp_0_13,tmp_0_14,tmp_0_15,tmp_0_16,tmp_0_17,tmp_0_18,tmp_0_19,tmp_0_20,tmp_0_21,tmp_0_22,tmp_0_23,tmp_0_24,tmp_0_25,tmp_0_26,tmp_0_27,tmp_0_28,tmp_0_29,tmp_0_30,tmp_0_31,tmp_0_32,tmp_0_33,tmp_0_34,tmp_0_35,tmp_0_36,tmp_0_37,tmp_0_38,tmp_0_39,tmp_0_40,tmp_0_41,tmp_0_42,tmp_0_43,tmp_0_44,tmp_0_45,tmp_0_46,tmp_0_47,tmp_0_48,tmp_0_49,tmp_0_50,tmp_0_51,tmp_0_52,tmp_0_53,tmp_0_54,tmp_0_55,tmp_0_56,tmp_0_57,tmp_0_58,tmp_0_59,tmp_0_60,tmp_0_61,tmp_0_62,tmp_0_63,tmp_0_64,tmp_0_65,tmp_0_66,tmp_0_67,tmp_0_68,tmp_0_69,tmp_0_70,tmp_0_71};
wire tmp_1_0;
assign tmp_1_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]);
wire tmp_1_1;
assign tmp_1_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]);
wire tmp_1_2;
assign tmp_1_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]);
wire tmp_1_3;
assign tmp_1_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]);
wire tmp_1_4;
assign tmp_1_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]);
wire tmp_1_5;
assign tmp_1_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]);
wire tmp_1_6;
assign tmp_1_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]);
wire tmp_1_7;
assign tmp_1_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]);
wire tmp_1_8;
assign tmp_1_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]);
wire tmp_1_9;
assign tmp_1_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]);
wire tmp_1_10;
assign tmp_1_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_1_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_1_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_1_V_read[10]);
wire tmp_1_11;
assign tmp_1_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]);
wire tmp_1_12;
assign tmp_1_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]);
wire tmp_1_14;
assign tmp_1_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]);
wire tmp_1_15;
assign tmp_1_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_1_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_1_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_1_V_read[15]);
wire tmp_1_16;
assign tmp_1_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]);
wire tmp_1_17;
assign tmp_1_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]);
wire tmp_1_18;
assign tmp_1_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]);
wire tmp_1_19;
assign tmp_1_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]);
wire tmp_1_20;
assign tmp_1_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]);
wire tmp_1_22;
assign tmp_1_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]);
wire tmp_1_23;
assign tmp_1_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_1_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_1_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_1_V_read[23]);
wire tmp_1_24;
assign tmp_1_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]);
wire tmp_1_25;
assign tmp_1_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]);
wire tmp_1_26;
assign tmp_1_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]);
wire tmp_1_27;
assign tmp_1_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]);
wire tmp_1_28;
assign tmp_1_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]);
wire tmp_1_30;
assign tmp_1_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]);
wire tmp_1_31;
assign tmp_1_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]);
wire tmp_1_32;
assign tmp_1_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]);
wire tmp_1_33;
assign tmp_1_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_1_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_1_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_1_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_1_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_1_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_1_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_1_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_1_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_1_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_1_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_1_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_1_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_1_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_1_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_1_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_1_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_1_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_1_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_1_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_1_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_1_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_1_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_1_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_1_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_1_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_1_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_1_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_1_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_1_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_1_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_1_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_1_V_read[33]);
wire tmp_1_34;
assign tmp_1_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_1_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_1_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_1_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_1_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_1_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_1_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_1_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_1_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_1_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_1_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_1_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_1_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_1_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_1_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_1_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_1_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_1_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_1_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_1_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_1_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_1_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_1_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_1_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_1_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_1_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_1_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_1_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_1_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_1_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_1_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_1_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_1_V_read[34]);
wire tmp_1_35;
assign tmp_1_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]);
wire tmp_1_36;
assign tmp_1_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]);
wire tmp_1_37;
assign tmp_1_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]);
wire tmp_1_38;
assign tmp_1_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]);
wire tmp_1_39;
assign tmp_1_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_1_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_1_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_1_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_1_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_1_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_1_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_1_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_1_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_1_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_1_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_1_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_1_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_1_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_1_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_1_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_1_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_1_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_1_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_1_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_1_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_1_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_1_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_1_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_1_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_1_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_1_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_1_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_1_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_1_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_1_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_1_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_1_V_read[39]);
wire tmp_1_40;
assign tmp_1_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]);
wire tmp_1_41;
assign tmp_1_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]);
wire tmp_1_42;
assign tmp_1_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]);
wire tmp_1_43;
assign tmp_1_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]);
wire tmp_1_44;
assign tmp_1_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]);
wire tmp_1_45;
assign tmp_1_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]);
wire tmp_1_46;
assign tmp_1_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]);
wire tmp_1_47;
assign tmp_1_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]);
wire tmp_1_48;
assign tmp_1_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]);
wire tmp_1_49;
assign tmp_1_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]);
wire tmp_1_50;
assign tmp_1_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]);
wire tmp_1_51;
assign tmp_1_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]);
wire tmp_1_52;
assign tmp_1_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]);
wire tmp_1_54;
assign tmp_1_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]);
wire tmp_1_55;
assign tmp_1_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_1_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_1_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_1_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_1_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_1_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_1_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_1_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_1_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_1_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_1_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_1_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_1_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_1_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_1_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_1_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_1_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_1_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_1_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_1_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_1_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_1_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_1_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_1_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_1_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_1_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_1_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_1_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_1_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_1_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_1_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_1_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_1_V_read[55]);
wire tmp_1_56;
assign tmp_1_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]);
wire tmp_1_57;
assign tmp_1_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]);
wire tmp_1_58;
assign tmp_1_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]);
wire tmp_1_59;
assign tmp_1_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]);
wire tmp_1_60;
assign tmp_1_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]);
wire tmp_1_61;
assign tmp_1_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]);
wire tmp_1_62;
assign tmp_1_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]);
wire tmp_1_63;
assign tmp_1_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]);
wire tmp_1_64;
assign tmp_1_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]);
wire tmp_1_65;
assign tmp_1_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]);
wire tmp_1_66;
assign tmp_1_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]);
wire tmp_1_67;
assign tmp_1_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]);
wire tmp_1_68;
assign tmp_1_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]);
wire tmp_1_69;
assign tmp_1_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]);
wire tmp_1_70;
assign tmp_1_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]);
wire tmp_1_71;
assign tmp_1_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]);
assign ap_return_1 = {tmp_1_0,tmp_1_1,tmp_1_2,tmp_1_3,tmp_1_4,tmp_1_5,tmp_1_6,tmp_1_7,tmp_1_8,tmp_1_9,tmp_1_10,tmp_1_11,tmp_1_12,1'b0,tmp_1_14,tmp_1_15,tmp_1_16,tmp_1_17,tmp_1_18,tmp_1_19,tmp_1_20,1'b0,tmp_1_22,tmp_1_23,tmp_1_24,tmp_1_25,tmp_1_26,tmp_1_27,tmp_1_28,1'b0,tmp_1_30,tmp_1_31,tmp_1_32,tmp_1_33,tmp_1_34,tmp_1_35,tmp_1_36,tmp_1_37,tmp_1_38,tmp_1_39,tmp_1_40,tmp_1_41,tmp_1_42,tmp_1_43,tmp_1_44,tmp_1_45,tmp_1_46,tmp_1_47,tmp_1_48,tmp_1_49,tmp_1_50,tmp_1_51,tmp_1_52,1'b0,tmp_1_54,tmp_1_55,tmp_1_56,tmp_1_57,tmp_1_58,tmp_1_59,tmp_1_60,tmp_1_61,tmp_1_62,tmp_1_63,tmp_1_64,tmp_1_65,tmp_1_66,tmp_1_67,tmp_1_68,tmp_1_69,tmp_1_70,tmp_1_71};
wire tmp_2_0;
assign tmp_2_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]);
wire tmp_2_1;
assign tmp_2_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]);
wire tmp_2_2;
assign tmp_2_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]);
wire tmp_2_3;
assign tmp_2_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]);
wire tmp_2_4;
assign tmp_2_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]);
wire tmp_2_5;
assign tmp_2_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]);
wire tmp_2_6;
assign tmp_2_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]);
wire tmp_2_7;
assign tmp_2_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]);
wire tmp_2_8;
assign tmp_2_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]);
wire tmp_2_9;
assign tmp_2_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]);
wire tmp_2_10;
assign tmp_2_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]);
wire tmp_2_11;
assign tmp_2_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]);
wire tmp_2_12;
assign tmp_2_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]);
wire tmp_2_14;
assign tmp_2_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_2_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_2_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_2_V_read[14]);
wire tmp_2_15;
assign tmp_2_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_2_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_2_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_2_V_read[15]);
wire tmp_2_16;
assign tmp_2_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]);
wire tmp_2_17;
assign tmp_2_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]);
wire tmp_2_18;
assign tmp_2_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]);
wire tmp_2_19;
assign tmp_2_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]);
wire tmp_2_20;
assign tmp_2_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]);
wire tmp_2_21;
assign tmp_2_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]);
wire tmp_2_22;
assign tmp_2_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]);
wire tmp_2_23;
assign tmp_2_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]);
wire tmp_2_24;
assign tmp_2_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]);
wire tmp_2_25;
assign tmp_2_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]);
wire tmp_2_26;
assign tmp_2_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]);
wire tmp_2_27;
assign tmp_2_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]);
wire tmp_2_28;
assign tmp_2_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_2_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_2_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_2_V_read[28]);
wire tmp_2_29;
assign tmp_2_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]);
wire tmp_2_30;
assign tmp_2_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]);
wire tmp_2_31;
assign tmp_2_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_2_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_2_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_2_V_read[31]);
wire tmp_2_32;
assign tmp_2_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]);
wire tmp_2_33;
assign tmp_2_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]);
wire tmp_2_34;
assign tmp_2_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]);
wire tmp_2_35;
assign tmp_2_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]);
wire tmp_2_36;
assign tmp_2_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]);
wire tmp_2_37;
assign tmp_2_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]);
wire tmp_2_38;
assign tmp_2_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]);
wire tmp_2_39;
assign tmp_2_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]);
wire tmp_2_40;
assign tmp_2_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]);
wire tmp_2_41;
assign tmp_2_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]);
wire tmp_2_42;
assign tmp_2_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]);
wire tmp_2_43;
assign tmp_2_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]);
wire tmp_2_44;
assign tmp_2_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]);
wire tmp_2_45;
assign tmp_2_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]);
wire tmp_2_46;
assign tmp_2_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]);
wire tmp_2_47;
assign tmp_2_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_2_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_2_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_2_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_2_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_2_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_2_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_2_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_2_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_2_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_2_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_2_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_2_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_2_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_2_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_2_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_2_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_2_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_2_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_2_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_2_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_2_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_2_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_2_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_2_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_2_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_2_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_2_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_2_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_2_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_2_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_2_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_2_V_read[47]);
wire tmp_2_48;
assign tmp_2_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]);
wire tmp_2_49;
assign tmp_2_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]);
wire tmp_2_50;
assign tmp_2_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]);
wire tmp_2_51;
assign tmp_2_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]);
wire tmp_2_52;
assign tmp_2_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]);
wire tmp_2_53;
assign tmp_2_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_2_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_2_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_2_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_2_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_2_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_2_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_2_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_2_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_2_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_2_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_2_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_2_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_2_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_2_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_2_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_2_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_2_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_2_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_2_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_2_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_2_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_2_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_2_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_2_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_2_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_2_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_2_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_2_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_2_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_2_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_2_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_2_V_read[53]);
wire tmp_2_54;
assign tmp_2_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]);
wire tmp_2_55;
assign tmp_2_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_2_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_2_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_2_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_2_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_2_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_2_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_2_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_2_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_2_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_2_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_2_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_2_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_2_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_2_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_2_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_2_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_2_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_2_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_2_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_2_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_2_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_2_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_2_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_2_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_2_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_2_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_2_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_2_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_2_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_2_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_2_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_2_V_read[55]);
wire tmp_2_56;
assign tmp_2_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]);
wire tmp_2_57;
assign tmp_2_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]);
wire tmp_2_58;
assign tmp_2_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_2_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_2_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_2_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_2_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_2_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_2_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_2_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_2_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_2_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_2_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_2_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_2_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_2_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_2_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_2_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_2_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_2_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_2_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_2_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_2_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_2_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_2_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_2_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_2_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_2_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_2_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_2_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_2_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_2_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_2_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_2_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_2_V_read[58]);
wire tmp_2_59;
assign tmp_2_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]);
wire tmp_2_60;
assign tmp_2_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]);
wire tmp_2_61;
assign tmp_2_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]);
wire tmp_2_62;
assign tmp_2_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]);
wire tmp_2_63;
assign tmp_2_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]);
wire tmp_2_64;
assign tmp_2_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_2_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_2_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_2_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_2_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_2_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_2_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_2_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_2_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_2_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_2_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_2_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_2_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_2_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_2_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_2_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_2_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_2_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_2_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_2_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_2_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_2_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_2_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_2_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_2_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_2_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_2_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_2_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_2_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_2_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_2_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_2_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_2_V_read[64]);
wire tmp_2_65;
assign tmp_2_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_2_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_2_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_2_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_2_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_2_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_2_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_2_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_2_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_2_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_2_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_2_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_2_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_2_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_2_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_2_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_2_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_2_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_2_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_2_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_2_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_2_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_2_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_2_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_2_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_2_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_2_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_2_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_2_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_2_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_2_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_2_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_2_V_read[65]);
wire tmp_2_66;
assign tmp_2_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]);
wire tmp_2_67;
assign tmp_2_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]);
wire tmp_2_68;
assign tmp_2_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]);
wire tmp_2_69;
assign tmp_2_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]);
wire tmp_2_70;
assign tmp_2_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]);
wire tmp_2_71;
assign tmp_2_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]);
assign ap_return_2 = {tmp_2_0,tmp_2_1,tmp_2_2,tmp_2_3,tmp_2_4,tmp_2_5,tmp_2_6,tmp_2_7,tmp_2_8,tmp_2_9,tmp_2_10,tmp_2_11,tmp_2_12,1'b0,tmp_2_14,tmp_2_15,tmp_2_16,tmp_2_17,tmp_2_18,tmp_2_19,tmp_2_20,tmp_2_21,tmp_2_22,tmp_2_23,tmp_2_24,tmp_2_25,tmp_2_26,tmp_2_27,tmp_2_28,tmp_2_29,tmp_2_30,tmp_2_31,tmp_2_32,tmp_2_33,tmp_2_34,tmp_2_35,tmp_2_36,tmp_2_37,tmp_2_38,tmp_2_39,tmp_2_40,tmp_2_41,tmp_2_42,tmp_2_43,tmp_2_44,tmp_2_45,tmp_2_46,tmp_2_47,tmp_2_48,tmp_2_49,tmp_2_50,tmp_2_51,tmp_2_52,tmp_2_53,tmp_2_54,tmp_2_55,tmp_2_56,tmp_2_57,tmp_2_58,tmp_2_59,tmp_2_60,tmp_2_61,tmp_2_62,tmp_2_63,tmp_2_64,tmp_2_65,tmp_2_66,tmp_2_67,tmp_2_68,tmp_2_69,tmp_2_70,tmp_2_71};
wire tmp_3_0;
assign tmp_3_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]);
wire tmp_3_1;
assign tmp_3_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]);
wire tmp_3_2;
assign tmp_3_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]);
wire tmp_3_3;
assign tmp_3_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]);
wire tmp_3_4;
assign tmp_3_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]);
wire tmp_3_5;
assign tmp_3_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]);
wire tmp_3_6;
assign tmp_3_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]);
wire tmp_3_7;
assign tmp_3_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]);
wire tmp_3_8;
assign tmp_3_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]);
wire tmp_3_9;
assign tmp_3_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]);
wire tmp_3_10;
assign tmp_3_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_3_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_3_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_3_V_read[10]);
wire tmp_3_11;
assign tmp_3_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]);
wire tmp_3_12;
assign tmp_3_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]);
wire tmp_3_13;
assign tmp_3_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]);
wire tmp_3_14;
assign tmp_3_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]);
wire tmp_3_15;
assign tmp_3_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_3_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_3_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_3_V_read[15]);
wire tmp_3_16;
assign tmp_3_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]);
wire tmp_3_17;
assign tmp_3_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]);
wire tmp_3_18;
assign tmp_3_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]);
wire tmp_3_19;
assign tmp_3_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]);
wire tmp_3_20;
assign tmp_3_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]);
wire tmp_3_21;
assign tmp_3_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]);
wire tmp_3_22;
assign tmp_3_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]);
wire tmp_3_23;
assign tmp_3_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]);
wire tmp_3_24;
assign tmp_3_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]);
wire tmp_3_25;
assign tmp_3_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]);
wire tmp_3_26;
assign tmp_3_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]);
wire tmp_3_27;
assign tmp_3_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]);
wire tmp_3_28;
assign tmp_3_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]);
wire tmp_3_29;
assign tmp_3_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]);
wire tmp_3_30;
assign tmp_3_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]);
wire tmp_3_31;
assign tmp_3_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_3_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_3_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_3_V_read[31]);
wire tmp_3_32;
assign tmp_3_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]);
wire tmp_3_33;
assign tmp_3_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]);
wire tmp_3_34;
assign tmp_3_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_3_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_3_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_3_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_3_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_3_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_3_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_3_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_3_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_3_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_3_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_3_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_3_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_3_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_3_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_3_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_3_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_3_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_3_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_3_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_3_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_3_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_3_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_3_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_3_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_3_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_3_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_3_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_3_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_3_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_3_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_3_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_3_V_read[34]);
wire tmp_3_35;
assign tmp_3_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]);
wire tmp_3_36;
assign tmp_3_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]);
wire tmp_3_37;
assign tmp_3_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_3_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_3_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_3_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_3_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_3_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_3_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_3_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_3_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_3_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_3_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_3_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_3_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_3_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_3_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_3_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_3_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_3_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_3_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_3_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_3_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_3_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_3_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_3_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_3_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_3_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_3_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_3_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_3_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_3_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_3_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_3_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_3_V_read[37]);
wire tmp_3_38;
assign tmp_3_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]);
wire tmp_3_39;
assign tmp_3_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_3_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_3_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_3_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_3_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_3_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_3_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_3_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_3_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_3_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_3_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_3_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_3_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_3_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_3_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_3_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_3_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_3_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_3_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_3_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_3_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_3_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_3_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_3_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_3_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_3_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_3_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_3_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_3_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_3_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_3_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_3_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_3_V_read[39]);
wire tmp_3_40;
assign tmp_3_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]);
wire tmp_3_41;
assign tmp_3_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]);
wire tmp_3_42;
assign tmp_3_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]);
wire tmp_3_43;
assign tmp_3_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_3_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_3_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_3_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_3_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_3_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_3_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_3_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_3_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_3_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_3_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_3_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_3_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_3_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_3_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_3_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_3_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_3_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_3_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_3_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_3_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_3_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_3_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_3_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_3_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_3_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_3_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_3_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_3_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_3_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_3_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_3_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_3_V_read[43]);
wire tmp_3_44;
assign tmp_3_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_3_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_3_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_3_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_3_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_3_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_3_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_3_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_3_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_3_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_3_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_3_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_3_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_3_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_3_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_3_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_3_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_3_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_3_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_3_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_3_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_3_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_3_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_3_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_3_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_3_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_3_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_3_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_3_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_3_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_3_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_3_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_3_V_read[44]);
wire tmp_3_45;
assign tmp_3_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]);
wire tmp_3_46;
assign tmp_3_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_3_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_3_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_3_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_3_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_3_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_3_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_3_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_3_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_3_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_3_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_3_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_3_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_3_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_3_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_3_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_3_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_3_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_3_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_3_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_3_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_3_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_3_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_3_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_3_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_3_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_3_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_3_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_3_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_3_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_3_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_3_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_3_V_read[46]);
wire tmp_3_47;
assign tmp_3_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_3_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_3_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_3_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_3_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_3_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_3_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_3_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_3_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_3_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_3_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_3_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_3_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_3_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_3_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_3_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_3_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_3_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_3_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_3_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_3_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_3_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_3_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_3_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_3_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_3_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_3_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_3_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_3_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_3_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_3_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_3_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_3_V_read[47]);
wire tmp_3_48;
assign tmp_3_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_3_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_3_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_3_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_3_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_3_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_3_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_3_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_3_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_3_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_3_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_3_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_3_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_3_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_3_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_3_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_3_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_3_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_3_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_3_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_3_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_3_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_3_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_3_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_3_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_3_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_3_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_3_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_3_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_3_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_3_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_3_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_3_V_read[48]);
wire tmp_3_49;
assign tmp_3_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]);
wire tmp_3_50;
assign tmp_3_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]);
wire tmp_3_51;
assign tmp_3_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]);
wire tmp_3_52;
assign tmp_3_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]);
wire tmp_3_53;
assign tmp_3_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]);
wire tmp_3_54;
assign tmp_3_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]);
wire tmp_3_55;
assign tmp_3_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]);
wire tmp_3_56;
assign tmp_3_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]);
wire tmp_3_57;
assign tmp_3_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]);
wire tmp_3_58;
assign tmp_3_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_3_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_3_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_3_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_3_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_3_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_3_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_3_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_3_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_3_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_3_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_3_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_3_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_3_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_3_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_3_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_3_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_3_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_3_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_3_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_3_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_3_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_3_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_3_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_3_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_3_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_3_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_3_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_3_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_3_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_3_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_3_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_3_V_read[58]);
wire tmp_3_59;
assign tmp_3_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]);
wire tmp_3_60;
assign tmp_3_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_3_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_3_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_3_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_3_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_3_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_3_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_3_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_3_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_3_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_3_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_3_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_3_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_3_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_3_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_3_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_3_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_3_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_3_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_3_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_3_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_3_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_3_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_3_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_3_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_3_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_3_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_3_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_3_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_3_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_3_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_3_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_3_V_read[60]);
wire tmp_3_61;
assign tmp_3_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]);
wire tmp_3_63;
assign tmp_3_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]);
wire tmp_3_64;
assign tmp_3_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_3_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_3_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_3_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_3_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_3_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_3_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_3_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_3_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_3_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_3_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_3_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_3_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_3_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_3_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_3_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_3_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_3_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_3_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_3_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_3_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_3_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_3_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_3_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_3_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_3_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_3_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_3_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_3_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_3_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_3_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_3_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_3_V_read[64]);
wire tmp_3_65;
assign tmp_3_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]);
wire tmp_3_66;
assign tmp_3_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]);
wire tmp_3_67;
assign tmp_3_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]);
wire tmp_3_68;
assign tmp_3_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]);
wire tmp_3_69;
assign tmp_3_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_3_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_3_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_3_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_3_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_3_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_3_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_3_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_3_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_3_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_3_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_3_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_3_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_3_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_3_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_3_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_3_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_3_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_3_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_3_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_3_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_3_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_3_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_3_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_3_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_3_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_3_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_3_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_3_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_3_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_3_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_3_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_3_V_read[69]);
wire tmp_3_70;
assign tmp_3_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]);
wire tmp_3_71;
assign tmp_3_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]);
assign ap_return_3 = {tmp_3_0,tmp_3_1,tmp_3_2,tmp_3_3,tmp_3_4,tmp_3_5,tmp_3_6,tmp_3_7,tmp_3_8,tmp_3_9,tmp_3_10,tmp_3_11,tmp_3_12,tmp_3_13,tmp_3_14,tmp_3_15,tmp_3_16,tmp_3_17,tmp_3_18,tmp_3_19,tmp_3_20,tmp_3_21,tmp_3_22,tmp_3_23,tmp_3_24,tmp_3_25,tmp_3_26,tmp_3_27,tmp_3_28,tmp_3_29,tmp_3_30,tmp_3_31,tmp_3_32,tmp_3_33,tmp_3_34,tmp_3_35,tmp_3_36,tmp_3_37,tmp_3_38,tmp_3_39,tmp_3_40,tmp_3_41,tmp_3_42,tmp_3_43,tmp_3_44,tmp_3_45,tmp_3_46,tmp_3_47,tmp_3_48,tmp_3_49,tmp_3_50,tmp_3_51,tmp_3_52,tmp_3_53,tmp_3_54,tmp_3_55,tmp_3_56,tmp_3_57,tmp_3_58,tmp_3_59,tmp_3_60,tmp_3_61,1'b0,tmp_3_63,tmp_3_64,tmp_3_65,tmp_3_66,tmp_3_67,tmp_3_68,tmp_3_69,tmp_3_70,tmp_3_71};
wire tmp_4_0;
assign tmp_4_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]);
wire tmp_4_1;
assign tmp_4_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]);
wire tmp_4_2;
assign tmp_4_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]);
wire tmp_4_3;
assign tmp_4_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]);
wire tmp_4_4;
assign tmp_4_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]);
wire tmp_4_6;
assign tmp_4_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]);
wire tmp_4_7;
assign tmp_4_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]);
wire tmp_4_8;
assign tmp_4_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]);
wire tmp_4_9;
assign tmp_4_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]);
wire tmp_4_10;
assign tmp_4_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_4_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_4_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_4_V_read[10]);
wire tmp_4_11;
assign tmp_4_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]);
wire tmp_4_12;
assign tmp_4_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]);
wire tmp_4_14;
assign tmp_4_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]);
wire tmp_4_15;
assign tmp_4_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_4_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_4_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_4_V_read[15]);
wire tmp_4_16;
assign tmp_4_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]);
wire tmp_4_17;
assign tmp_4_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]);
wire tmp_4_18;
assign tmp_4_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]);
wire tmp_4_19;
assign tmp_4_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]);
wire tmp_4_20;
assign tmp_4_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]);
wire tmp_4_21;
assign tmp_4_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]);
wire tmp_4_22;
assign tmp_4_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]);
wire tmp_4_23;
assign tmp_4_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]);
wire tmp_4_24;
assign tmp_4_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]);
wire tmp_4_25;
assign tmp_4_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_4_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_4_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_4_V_read[25]);
wire tmp_4_26;
assign tmp_4_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]);
wire tmp_4_27;
assign tmp_4_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]);
wire tmp_4_28;
assign tmp_4_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]);
wire tmp_4_30;
assign tmp_4_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]);
wire tmp_4_31;
assign tmp_4_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]);
wire tmp_4_32;
assign tmp_4_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]);
wire tmp_4_33;
assign tmp_4_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]);
wire tmp_4_34;
assign tmp_4_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]);
wire tmp_4_35;
assign tmp_4_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]);
wire tmp_4_36;
assign tmp_4_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]);
wire tmp_4_37;
assign tmp_4_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]);
wire tmp_4_38;
assign tmp_4_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]);
wire tmp_4_39;
assign tmp_4_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]);
wire tmp_4_40;
assign tmp_4_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]);
wire tmp_4_41;
assign tmp_4_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]);
wire tmp_4_42;
assign tmp_4_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]);
wire tmp_4_43;
assign tmp_4_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]);
wire tmp_4_44;
assign tmp_4_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]);
wire tmp_4_45;
assign tmp_4_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]);
wire tmp_4_46;
assign tmp_4_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_4_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_4_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_4_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_4_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_4_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_4_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_4_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_4_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_4_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_4_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_4_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_4_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_4_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_4_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_4_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_4_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_4_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_4_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_4_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_4_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_4_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_4_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_4_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_4_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_4_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_4_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_4_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_4_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_4_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_4_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_4_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_4_V_read[46]);
wire tmp_4_47;
assign tmp_4_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]);
wire tmp_4_48;
assign tmp_4_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]);
wire tmp_4_49;
assign tmp_4_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]);
wire tmp_4_50;
assign tmp_4_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]);
wire tmp_4_51;
assign tmp_4_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]);
wire tmp_4_52;
assign tmp_4_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]);
wire tmp_4_53;
assign tmp_4_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]);
wire tmp_4_54;
assign tmp_4_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]);
wire tmp_4_55;
assign tmp_4_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]);
wire tmp_4_56;
assign tmp_4_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]);
wire tmp_4_57;
assign tmp_4_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]);
wire tmp_4_58;
assign tmp_4_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]);
wire tmp_4_59;
assign tmp_4_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]);
wire tmp_4_60;
assign tmp_4_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]);
wire tmp_4_62;
assign tmp_4_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_4_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_4_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_4_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_4_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_4_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_4_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_4_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_4_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_4_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_4_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_4_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_4_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_4_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_4_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_4_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_4_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_4_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_4_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_4_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_4_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_4_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_4_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_4_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_4_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_4_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_4_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_4_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_4_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_4_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_4_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_4_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_4_V_read[62]);
wire tmp_4_63;
assign tmp_4_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]);
wire tmp_4_64;
assign tmp_4_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]);
wire tmp_4_65;
assign tmp_4_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]);
wire tmp_4_66;
assign tmp_4_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]);
wire tmp_4_67;
assign tmp_4_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]);
wire tmp_4_68;
assign tmp_4_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]);
wire tmp_4_70;
assign tmp_4_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]);
wire tmp_4_71;
assign tmp_4_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_4_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_4_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_4_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_4_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_4_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_4_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_4_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_4_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_4_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_4_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_4_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_4_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_4_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_4_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_4_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_4_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_4_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_4_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_4_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_4_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_4_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_4_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_4_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_4_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_4_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_4_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_4_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_4_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_4_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_4_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_4_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_4_V_read[71]);
assign ap_return_4 = {tmp_4_0,tmp_4_1,tmp_4_2,tmp_4_3,tmp_4_4,1'b0,tmp_4_6,tmp_4_7,tmp_4_8,tmp_4_9,tmp_4_10,tmp_4_11,tmp_4_12,1'b0,tmp_4_14,tmp_4_15,tmp_4_16,tmp_4_17,tmp_4_18,tmp_4_19,tmp_4_20,tmp_4_21,tmp_4_22,tmp_4_23,tmp_4_24,tmp_4_25,tmp_4_26,tmp_4_27,tmp_4_28,1'b0,tmp_4_30,tmp_4_31,tmp_4_32,tmp_4_33,tmp_4_34,tmp_4_35,tmp_4_36,tmp_4_37,tmp_4_38,tmp_4_39,tmp_4_40,tmp_4_41,tmp_4_42,tmp_4_43,tmp_4_44,tmp_4_45,tmp_4_46,tmp_4_47,tmp_4_48,tmp_4_49,tmp_4_50,tmp_4_51,tmp_4_52,tmp_4_53,tmp_4_54,tmp_4_55,tmp_4_56,tmp_4_57,tmp_4_58,tmp_4_59,tmp_4_60,1'b0,tmp_4_62,tmp_4_63,tmp_4_64,tmp_4_65,tmp_4_66,tmp_4_67,tmp_4_68,1'b0,tmp_4_70,tmp_4_71};
wire tmp_5_0;
assign tmp_5_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]);
wire tmp_5_1;
assign tmp_5_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]);
wire tmp_5_2;
assign tmp_5_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]);
wire tmp_5_3;
assign tmp_5_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]);
wire tmp_5_4;
assign tmp_5_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]);
wire tmp_5_6;
assign tmp_5_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]);
wire tmp_5_7;
assign tmp_5_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]);
wire tmp_5_8;
assign tmp_5_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]);
wire tmp_5_9;
assign tmp_5_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]);
wire tmp_5_10;
assign tmp_5_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]);
wire tmp_5_11;
assign tmp_5_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]);
wire tmp_5_12;
assign tmp_5_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]);
wire tmp_5_13;
assign tmp_5_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]);
wire tmp_5_14;
assign tmp_5_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_5_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_5_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_5_V_read[14]);
wire tmp_5_15;
assign tmp_5_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_5_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_5_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_5_V_read[15]);
wire tmp_5_16;
assign tmp_5_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]);
wire tmp_5_17;
assign tmp_5_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]);
wire tmp_5_18;
assign tmp_5_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]);
wire tmp_5_19;
assign tmp_5_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]);
wire tmp_5_20;
assign tmp_5_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]);
wire tmp_5_21;
assign tmp_5_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]);
wire tmp_5_22;
assign tmp_5_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]);
wire tmp_5_23;
assign tmp_5_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]);
wire tmp_5_24;
assign tmp_5_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]);
wire tmp_5_25;
assign tmp_5_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]);
wire tmp_5_26;
assign tmp_5_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]);
wire tmp_5_27;
assign tmp_5_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]);
wire tmp_5_28;
assign tmp_5_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]);
wire tmp_5_29;
assign tmp_5_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]);
wire tmp_5_30;
assign tmp_5_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]);
wire tmp_5_31;
assign tmp_5_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]);
wire tmp_5_32;
assign tmp_5_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]);
wire tmp_5_33;
assign tmp_5_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]);
wire tmp_5_34;
assign tmp_5_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_5_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_5_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_5_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_5_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_5_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_5_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_5_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_5_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_5_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_5_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_5_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_5_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_5_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_5_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_5_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_5_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_5_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_5_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_5_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_5_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_5_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_5_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_5_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_5_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_5_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_5_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_5_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_5_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_5_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_5_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_5_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_5_V_read[34]);
wire tmp_5_35;
assign tmp_5_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]);
wire tmp_5_36;
assign tmp_5_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]);
wire tmp_5_37;
assign tmp_5_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]);
wire tmp_5_38;
assign tmp_5_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]);
wire tmp_5_39;
assign tmp_5_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_5_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_5_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_5_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_5_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_5_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_5_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_5_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_5_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_5_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_5_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_5_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_5_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_5_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_5_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_5_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_5_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_5_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_5_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_5_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_5_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_5_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_5_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_5_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_5_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_5_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_5_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_5_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_5_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_5_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_5_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_5_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_5_V_read[39]);
wire tmp_5_40;
assign tmp_5_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]);
wire tmp_5_41;
assign tmp_5_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]);
wire tmp_5_42;
assign tmp_5_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]);
wire tmp_5_43;
assign tmp_5_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]);
wire tmp_5_44;
assign tmp_5_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]);
wire tmp_5_45;
assign tmp_5_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]);
wire tmp_5_46;
assign tmp_5_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_5_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_5_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_5_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_5_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_5_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_5_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_5_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_5_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_5_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_5_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_5_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_5_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_5_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_5_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_5_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_5_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_5_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_5_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_5_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_5_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_5_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_5_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_5_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_5_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_5_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_5_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_5_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_5_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_5_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_5_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_5_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_5_V_read[46]);
wire tmp_5_47;
assign tmp_5_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]);
wire tmp_5_48;
assign tmp_5_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]);
wire tmp_5_49;
assign tmp_5_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]);
wire tmp_5_50;
assign tmp_5_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]);
wire tmp_5_51;
assign tmp_5_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]);
wire tmp_5_52;
assign tmp_5_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]);
wire tmp_5_53;
assign tmp_5_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]);
wire tmp_5_54;
assign tmp_5_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]);
wire tmp_5_55;
assign tmp_5_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]);
wire tmp_5_56;
assign tmp_5_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]);
wire tmp_5_57;
assign tmp_5_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]);
wire tmp_5_58;
assign tmp_5_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_5_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_5_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_5_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_5_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_5_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_5_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_5_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_5_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_5_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_5_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_5_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_5_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_5_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_5_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_5_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_5_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_5_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_5_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_5_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_5_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_5_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_5_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_5_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_5_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_5_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_5_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_5_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_5_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_5_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_5_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_5_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_5_V_read[58]);
wire tmp_5_59;
assign tmp_5_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]);
wire tmp_5_60;
assign tmp_5_60 = (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]);
wire tmp_5_61;
assign tmp_5_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]);
wire tmp_5_62;
assign tmp_5_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]);
wire tmp_5_63;
assign tmp_5_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]);
wire tmp_5_64;
assign tmp_5_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]);
wire tmp_5_65;
assign tmp_5_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]);
wire tmp_5_66;
assign tmp_5_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]);
wire tmp_5_67;
assign tmp_5_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]);
wire tmp_5_68;
assign tmp_5_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]);
wire tmp_5_69;
assign tmp_5_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]);
wire tmp_5_70;
assign tmp_5_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]);
wire tmp_5_71;
assign tmp_5_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]);
assign ap_return_5 = {tmp_5_0,tmp_5_1,tmp_5_2,tmp_5_3,tmp_5_4,1'b0,tmp_5_6,tmp_5_7,tmp_5_8,tmp_5_9,tmp_5_10,tmp_5_11,tmp_5_12,tmp_5_13,tmp_5_14,tmp_5_15,tmp_5_16,tmp_5_17,tmp_5_18,tmp_5_19,tmp_5_20,tmp_5_21,tmp_5_22,tmp_5_23,tmp_5_24,tmp_5_25,tmp_5_26,tmp_5_27,tmp_5_28,tmp_5_29,tmp_5_30,tmp_5_31,tmp_5_32,tmp_5_33,tmp_5_34,tmp_5_35,tmp_5_36,tmp_5_37,tmp_5_38,tmp_5_39,tmp_5_40,tmp_5_41,tmp_5_42,tmp_5_43,tmp_5_44,tmp_5_45,tmp_5_46,tmp_5_47,tmp_5_48,tmp_5_49,tmp_5_50,tmp_5_51,tmp_5_52,tmp_5_53,tmp_5_54,tmp_5_55,tmp_5_56,tmp_5_57,tmp_5_58,tmp_5_59,tmp_5_60,tmp_5_61,tmp_5_62,tmp_5_63,tmp_5_64,tmp_5_65,tmp_5_66,tmp_5_67,tmp_5_68,tmp_5_69,tmp_5_70,tmp_5_71};
wire tmp_6_0;
assign tmp_6_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]);
wire tmp_6_1;
assign tmp_6_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]);
wire tmp_6_2;
assign tmp_6_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]);
wire tmp_6_3;
assign tmp_6_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]);
wire tmp_6_4;
assign tmp_6_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]);
wire tmp_6_5;
assign tmp_6_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]);
wire tmp_6_6;
assign tmp_6_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]);
wire tmp_6_7;
assign tmp_6_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_6_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_6_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_6_V_read[7]);
wire tmp_6_8;
assign tmp_6_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_6_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_6_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_6_V_read[8]);
wire tmp_6_9;
assign tmp_6_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]);
wire tmp_6_10;
assign tmp_6_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]);
wire tmp_6_11;
assign tmp_6_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]);
wire tmp_6_12;
assign tmp_6_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]);
wire tmp_6_14;
assign tmp_6_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]);
wire tmp_6_15;
assign tmp_6_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]);
wire tmp_6_16;
assign tmp_6_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]);
wire tmp_6_17;
assign tmp_6_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]);
wire tmp_6_18;
assign tmp_6_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]);
wire tmp_6_19;
assign tmp_6_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]);
wire tmp_6_20;
assign tmp_6_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]);
wire tmp_6_21;
assign tmp_6_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]);
wire tmp_6_22;
assign tmp_6_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]);
wire tmp_6_23;
assign tmp_6_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_6_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_6_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_6_V_read[23]);
wire tmp_6_24;
assign tmp_6_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]);
wire tmp_6_25;
assign tmp_6_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]);
wire tmp_6_26;
assign tmp_6_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]);
wire tmp_6_27;
assign tmp_6_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]);
wire tmp_6_28;
assign tmp_6_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]);
wire tmp_6_29;
assign tmp_6_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]);
wire tmp_6_30;
assign tmp_6_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]);
wire tmp_6_31;
assign tmp_6_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]);
wire tmp_6_32;
assign tmp_6_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]);
wire tmp_6_33;
assign tmp_6_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]);
wire tmp_6_34;
assign tmp_6_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_6_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_6_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_6_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_6_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_6_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_6_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_6_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_6_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_6_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_6_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_6_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_6_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_6_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_6_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_6_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_6_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_6_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_6_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_6_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_6_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_6_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_6_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_6_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_6_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_6_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_6_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_6_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_6_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_6_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_6_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_6_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_6_V_read[34]);
wire tmp_6_35;
assign tmp_6_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_6_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_6_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_6_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_6_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_6_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_6_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_6_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_6_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_6_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_6_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_6_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_6_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_6_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_6_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_6_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_6_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_6_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_6_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_6_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_6_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_6_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_6_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_6_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_6_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_6_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_6_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_6_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_6_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_6_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_6_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_6_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_6_V_read[35]);
wire tmp_6_36;
assign tmp_6_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]);
wire tmp_6_37;
assign tmp_6_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]);
wire tmp_6_38;
assign tmp_6_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]);
wire tmp_6_39;
assign tmp_6_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]);
wire tmp_6_40;
assign tmp_6_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]);
wire tmp_6_41;
assign tmp_6_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]);
wire tmp_6_42;
assign tmp_6_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]);
wire tmp_6_43;
assign tmp_6_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]);
wire tmp_6_44;
assign tmp_6_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]);
wire tmp_6_45;
assign tmp_6_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]);
wire tmp_6_46;
assign tmp_6_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]);
wire tmp_6_47;
assign tmp_6_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]);
wire tmp_6_48;
assign tmp_6_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]);
wire tmp_6_49;
assign tmp_6_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]);
wire tmp_6_50;
assign tmp_6_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]);
wire tmp_6_51;
assign tmp_6_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]);
wire tmp_6_52;
assign tmp_6_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]);
wire tmp_6_53;
assign tmp_6_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]);
wire tmp_6_54;
assign tmp_6_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_6_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_6_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_6_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_6_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_6_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_6_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_6_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_6_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_6_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_6_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_6_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_6_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_6_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_6_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_6_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_6_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_6_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_6_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_6_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_6_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_6_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_6_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_6_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_6_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_6_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_6_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_6_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_6_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_6_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_6_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_6_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_6_V_read[54]);
wire tmp_6_55;
assign tmp_6_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]);
wire tmp_6_56;
assign tmp_6_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]);
wire tmp_6_57;
assign tmp_6_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]);
wire tmp_6_58;
assign tmp_6_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]);
wire tmp_6_59;
assign tmp_6_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]);
wire tmp_6_60;
assign tmp_6_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]);
wire tmp_6_61;
assign tmp_6_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]);
wire tmp_6_62;
assign tmp_6_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_6_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_6_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_6_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_6_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_6_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_6_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_6_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_6_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_6_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_6_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_6_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_6_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_6_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_6_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_6_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_6_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_6_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_6_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_6_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_6_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_6_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_6_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_6_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_6_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_6_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_6_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_6_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_6_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_6_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_6_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_6_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_6_V_read[62]);
wire tmp_6_63;
assign tmp_6_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]);
wire tmp_6_64;
assign tmp_6_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]);
wire tmp_6_65;
assign tmp_6_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]);
wire tmp_6_66;
assign tmp_6_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]);
wire tmp_6_67;
assign tmp_6_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]);
wire tmp_6_68;
assign tmp_6_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]);
wire tmp_6_69;
assign tmp_6_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]);
wire tmp_6_70;
assign tmp_6_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]);
wire tmp_6_71;
assign tmp_6_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]);
assign ap_return_6 = {tmp_6_0,tmp_6_1,tmp_6_2,tmp_6_3,tmp_6_4,tmp_6_5,tmp_6_6,tmp_6_7,tmp_6_8,tmp_6_9,tmp_6_10,tmp_6_11,tmp_6_12,1'b0,tmp_6_14,tmp_6_15,tmp_6_16,tmp_6_17,tmp_6_18,tmp_6_19,tmp_6_20,tmp_6_21,tmp_6_22,tmp_6_23,tmp_6_24,tmp_6_25,tmp_6_26,tmp_6_27,tmp_6_28,tmp_6_29,tmp_6_30,tmp_6_31,tmp_6_32,tmp_6_33,tmp_6_34,tmp_6_35,tmp_6_36,tmp_6_37,tmp_6_38,tmp_6_39,tmp_6_40,tmp_6_41,tmp_6_42,tmp_6_43,tmp_6_44,tmp_6_45,tmp_6_46,tmp_6_47,tmp_6_48,tmp_6_49,tmp_6_50,tmp_6_51,tmp_6_52,tmp_6_53,tmp_6_54,tmp_6_55,tmp_6_56,tmp_6_57,tmp_6_58,tmp_6_59,tmp_6_60,tmp_6_61,tmp_6_62,tmp_6_63,tmp_6_64,tmp_6_65,tmp_6_66,tmp_6_67,tmp_6_68,tmp_6_69,tmp_6_70,tmp_6_71};
wire tmp_7_0;
assign tmp_7_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]);
wire tmp_7_1;
assign tmp_7_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]);
wire tmp_7_2;
assign tmp_7_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]);
wire tmp_7_3;
assign tmp_7_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]);
wire tmp_7_4;
assign tmp_7_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]);
wire tmp_7_5;
assign tmp_7_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]);
wire tmp_7_6;
assign tmp_7_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]);
wire tmp_7_7;
assign tmp_7_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]);
wire tmp_7_8;
assign tmp_7_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_7_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_7_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_7_V_read[8]);
wire tmp_7_9;
assign tmp_7_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]);
wire tmp_7_10;
assign tmp_7_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]);
wire tmp_7_11;
assign tmp_7_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_7_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_7_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_7_V_read[11]);
wire tmp_7_12;
assign tmp_7_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]);
wire tmp_7_13;
assign tmp_7_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]);
wire tmp_7_14;
assign tmp_7_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]);
wire tmp_7_15;
assign tmp_7_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]);
wire tmp_7_16;
assign tmp_7_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]);
wire tmp_7_17;
assign tmp_7_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]);
wire tmp_7_18;
assign tmp_7_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]);
wire tmp_7_19;
assign tmp_7_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]);
wire tmp_7_20;
assign tmp_7_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]);
wire tmp_7_21;
assign tmp_7_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]);
wire tmp_7_22;
assign tmp_7_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]);
wire tmp_7_23;
assign tmp_7_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]);
wire tmp_7_24;
assign tmp_7_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]);
wire tmp_7_25;
assign tmp_7_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_7_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_7_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_7_V_read[25]);
wire tmp_7_26;
assign tmp_7_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]);
wire tmp_7_27;
assign tmp_7_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]);
wire tmp_7_28;
assign tmp_7_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]);
wire tmp_7_30;
assign tmp_7_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]);
wire tmp_7_31;
assign tmp_7_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]);
wire tmp_7_32;
assign tmp_7_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]);
wire tmp_7_33;
assign tmp_7_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]);
wire tmp_7_34;
assign tmp_7_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]);
wire tmp_7_35;
assign tmp_7_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]);
wire tmp_7_36;
assign tmp_7_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]);
wire tmp_7_38;
assign tmp_7_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]);
wire tmp_7_39;
assign tmp_7_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_7_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_7_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_7_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_7_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_7_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_7_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_7_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_7_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_7_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_7_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_7_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_7_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_7_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_7_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_7_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_7_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_7_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_7_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_7_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_7_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_7_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_7_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_7_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_7_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_7_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_7_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_7_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_7_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_7_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_7_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_7_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_7_V_read[39]);
wire tmp_7_40;
assign tmp_7_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]);
wire tmp_7_41;
assign tmp_7_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]);
wire tmp_7_42;
assign tmp_7_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]);
wire tmp_7_43;
assign tmp_7_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]);
wire tmp_7_44;
assign tmp_7_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]);
wire tmp_7_45;
assign tmp_7_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]);
wire tmp_7_46;
assign tmp_7_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]);
wire tmp_7_47;
assign tmp_7_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]);
wire tmp_7_48;
assign tmp_7_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]);
wire tmp_7_49;
assign tmp_7_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]);
wire tmp_7_50;
assign tmp_7_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]);
wire tmp_7_51;
assign tmp_7_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]);
wire tmp_7_52;
assign tmp_7_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]);
wire tmp_7_54;
assign tmp_7_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]);
wire tmp_7_55;
assign tmp_7_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]);
wire tmp_7_56;
assign tmp_7_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]);
wire tmp_7_57;
assign tmp_7_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]);
wire tmp_7_58;
assign tmp_7_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]);
wire tmp_7_59;
assign tmp_7_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_7_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_7_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_7_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_7_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_7_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_7_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_7_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_7_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_7_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_7_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_7_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_7_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_7_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_7_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_7_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_7_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_7_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_7_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_7_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_7_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_7_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_7_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_7_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_7_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_7_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_7_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_7_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_7_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_7_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_7_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_7_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_7_V_read[59]);
wire tmp_7_60;
assign tmp_7_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]);
wire tmp_7_61;
assign tmp_7_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]);
wire tmp_7_62;
assign tmp_7_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]);
wire tmp_7_63;
assign tmp_7_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_7_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_7_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_7_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_7_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_7_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_7_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_7_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_7_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_7_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_7_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_7_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_7_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_7_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_7_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_7_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_7_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_7_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_7_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_7_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_7_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_7_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_7_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_7_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_7_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_7_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_7_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_7_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_7_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_7_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_7_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_7_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_7_V_read[63]);
wire tmp_7_64;
assign tmp_7_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]);
wire tmp_7_65;
assign tmp_7_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]);
wire tmp_7_66;
assign tmp_7_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]);
wire tmp_7_67;
assign tmp_7_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]);
wire tmp_7_68;
assign tmp_7_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]);
wire tmp_7_69;
assign tmp_7_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]);
wire tmp_7_70;
assign tmp_7_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]);
wire tmp_7_71;
assign tmp_7_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_7_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_7_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_7_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_7_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_7_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_7_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_7_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_7_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_7_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_7_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_7_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_7_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_7_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_7_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_7_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_7_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_7_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_7_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_7_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_7_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_7_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_7_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_7_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_7_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_7_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_7_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_7_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_7_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_7_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_7_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_7_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_7_V_read[71]);
assign ap_return_7 = {tmp_7_0,tmp_7_1,tmp_7_2,tmp_7_3,tmp_7_4,tmp_7_5,tmp_7_6,tmp_7_7,tmp_7_8,tmp_7_9,tmp_7_10,tmp_7_11,tmp_7_12,tmp_7_13,tmp_7_14,tmp_7_15,tmp_7_16,tmp_7_17,tmp_7_18,tmp_7_19,tmp_7_20,tmp_7_21,tmp_7_22,tmp_7_23,tmp_7_24,tmp_7_25,tmp_7_26,tmp_7_27,tmp_7_28,1'b0,tmp_7_30,tmp_7_31,tmp_7_32,tmp_7_33,tmp_7_34,tmp_7_35,tmp_7_36,1'b0,tmp_7_38,tmp_7_39,tmp_7_40,tmp_7_41,tmp_7_42,tmp_7_43,tmp_7_44,tmp_7_45,tmp_7_46,tmp_7_47,tmp_7_48,tmp_7_49,tmp_7_50,tmp_7_51,tmp_7_52,1'b0,tmp_7_54,tmp_7_55,tmp_7_56,tmp_7_57,tmp_7_58,tmp_7_59,tmp_7_60,tmp_7_61,tmp_7_62,tmp_7_63,tmp_7_64,tmp_7_65,tmp_7_66,tmp_7_67,tmp_7_68,tmp_7_69,tmp_7_70,tmp_7_71};
endmodule