`timescale 1 ns / 1 ps

module LUTARRAY_36u_8u_s (
        in_V,
        in_1_V,
        in_2_V,
        in_3_V,
        weight_0_0_V_read,
        weight_0_1_V_read,
        weight_0_2_V_read,
        weight_0_3_V_read,
        weight_0_4_V_read,
        weight_0_5_V_read,
        weight_0_6_V_read,
        weight_0_7_V_read,
        weight_0_8_V_read,
        weight_0_9_V_read,
        weight_0_10_V_read,
        weight_0_11_V_read,
        weight_0_12_V_read,
        weight_0_13_V_read,
        weight_0_14_V_read,
        weight_0_15_V_read,
        ap_return_0,
        ap_return_1,
        ap_return_2,
        ap_return_3,
        ap_return_4,
        ap_return_5,
        ap_return_6,
        ap_return_7,
        ap_return_8,
        ap_return_9,
        ap_return_10,
        ap_return_11,
        ap_return_12,
        ap_return_13,
        ap_return_14,
        ap_return_15);



input  [71:0] in_V;
input  [71:0] in_1_V;
input  [71:0] in_2_V;
input  [71:0] in_3_V;
input  [95:0] weight_0_0_V_read;
input  [95:0] weight_0_1_V_read;
input  [95:0] weight_0_2_V_read;
input  [95:0] weight_0_3_V_read;
input  [95:0] weight_0_4_V_read;
input  [95:0] weight_0_5_V_read;
input  [95:0] weight_0_6_V_read;
input  [95:0] weight_0_7_V_read;
input  [95:0] weight_0_8_V_read;
input  [95:0] weight_0_9_V_read;
input  [95:0] weight_0_10_V_read;
input  [95:0] weight_0_11_V_read;
input  [95:0] weight_0_12_V_read;
input  [95:0] weight_0_13_V_read;
input  [95:0] weight_0_14_V_read;
input  [95:0] weight_0_15_V_read;
output  [71:0] ap_return_0;
output  [71:0] ap_return_1;
output  [71:0] ap_return_2;
output  [71:0] ap_return_3;
output  [71:0] ap_return_4;
output  [71:0] ap_return_5;
output  [71:0] ap_return_6;
output  [71:0] ap_return_7;
output  [71:0] ap_return_8;
output  [71:0] ap_return_9;
output  [71:0] ap_return_10;
output  [71:0] ap_return_11;
output  [71:0] ap_return_12;
output  [71:0] ap_return_13;
output  [71:0] ap_return_14;
output  [71:0] ap_return_15;
wire tmp_0_1;
assign tmp_0_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_0_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_0_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_0_V_read[1]);
wire tmp_0_2;
assign tmp_0_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_0_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_0_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_0_V_read[2]);
wire tmp_0_3;
assign tmp_0_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_0_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_0_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_0_V_read[3]);
wire tmp_0_4;
assign tmp_0_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_0_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_0_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_0_V_read[4]);
wire tmp_0_5;
assign tmp_0_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_0_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_0_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_0_V_read[5]);
wire tmp_0_6;
assign tmp_0_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_0_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_0_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_0_V_read[6]);
wire tmp_0_8;
assign tmp_0_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_0_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_0_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_0_V_read[8]);
wire tmp_0_10;
assign tmp_0_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_0_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_0_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_0_V_read[10]);
wire tmp_0_11;
assign tmp_0_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_0_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_0_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_0_V_read[11]);
wire tmp_0_12;
assign tmp_0_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_0_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_0_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_0_V_read[12]);
wire tmp_0_13;
assign tmp_0_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_0_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_0_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_0_V_read[13]);
wire tmp_0_14;
assign tmp_0_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_0_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_0_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_0_V_read[14]);
wire tmp_0_15;
assign tmp_0_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_0_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_0_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_0_V_read[15]);
wire tmp_0_16;
assign tmp_0_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_0_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_0_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_0_V_read[16]);
wire tmp_0_17;
assign tmp_0_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_0_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_0_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_0_V_read[17]);
wire tmp_0_18;
assign tmp_0_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_0_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_0_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_0_V_read[18]);
wire tmp_0_19;
assign tmp_0_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_0_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_0_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_0_V_read[19]);
wire tmp_0_20;
assign tmp_0_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_0_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_0_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_0_V_read[20]);
wire tmp_0_21;
assign tmp_0_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_0_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_0_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_0_V_read[21]);
wire tmp_0_22;
assign tmp_0_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_0_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_0_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_0_V_read[22]);
wire tmp_0_23;
assign tmp_0_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_0_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_0_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_0_V_read[23]);
wire tmp_0_24;
assign tmp_0_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_0_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_0_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_0_V_read[24]);
wire tmp_0_25;
assign tmp_0_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_0_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_0_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_0_V_read[25]);
wire tmp_0_27;
assign tmp_0_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_0_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_0_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_0_V_read[27]);
wire tmp_0_28;
assign tmp_0_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_0_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_0_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_0_V_read[28]);
wire tmp_0_30;
assign tmp_0_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_0_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_0_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_0_V_read[30]);
wire tmp_0_32;
assign tmp_0_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_0_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_0_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_0_V_read[32]);
wire tmp_0_33;
assign tmp_0_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_0_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_0_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_0_V_read[33]);
wire tmp_0_34;
assign tmp_0_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_0_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_0_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_0_V_read[34]);
wire tmp_0_35;
assign tmp_0_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_0_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_0_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_0_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_0_V_read[35]);
wire tmp_0_36;
assign tmp_0_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_0_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_0_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_0_V_read[36]);
wire tmp_0_37;
assign tmp_0_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_0_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_0_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_0_V_read[37]);
wire tmp_0_40;
assign tmp_0_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_0_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_0_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_0_V_read[40]);
wire tmp_0_41;
assign tmp_0_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_0_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_0_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_0_V_read[41]);
wire tmp_0_42;
assign tmp_0_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_0_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_0_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_0_V_read[42]);
wire tmp_0_43;
assign tmp_0_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_0_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_0_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_0_V_read[43]);
wire tmp_0_44;
assign tmp_0_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_0_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_0_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_0_V_read[44]);
wire tmp_0_45;
assign tmp_0_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_0_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_0_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_0_V_read[45]);
wire tmp_0_46;
assign tmp_0_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_0_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_0_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_0_V_read[46]);
wire tmp_0_48;
assign tmp_0_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_0_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_0_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_0_V_read[48]);
wire tmp_0_49;
assign tmp_0_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_0_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_0_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_0_V_read[49]);
wire tmp_0_50;
assign tmp_0_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_0_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_0_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_0_V_read[50]);
wire tmp_0_51;
assign tmp_0_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_0_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_0_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_0_V_read[51]);
wire tmp_0_52;
assign tmp_0_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_0_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_0_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_0_V_read[52]);
wire tmp_0_53;
assign tmp_0_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_0_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_0_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_0_V_read[53]);
wire tmp_0_54;
assign tmp_0_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_0_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_0_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_0_V_read[54]);
wire tmp_0_55;
assign tmp_0_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_0_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_0_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_0_V_read[55]);
wire tmp_0_56;
assign tmp_0_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_0_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_0_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_0_V_read[56]);
wire tmp_0_57;
assign tmp_0_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_0_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_0_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_0_V_read[57]);
wire tmp_0_58;
assign tmp_0_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_0_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_0_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_0_V_read[58]);
wire tmp_0_59;
assign tmp_0_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_0_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_0_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_0_V_read[59]);
wire tmp_0_60;
assign tmp_0_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_0_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_0_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_0_V_read[60]);
wire tmp_0_61;
assign tmp_0_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_0_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_0_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_0_V_read[61]);
wire tmp_0_62;
assign tmp_0_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_0_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_0_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_0_V_read[62]);
wire tmp_0_63;
assign tmp_0_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_0_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_0_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_0_V_read[63]);
wire tmp_0_64;
assign tmp_0_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_0_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_0_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_0_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_0_V_read[64]);
wire tmp_0_65;
assign tmp_0_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_0_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_0_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_0_V_read[65]);
wire tmp_0_66;
assign tmp_0_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_0_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_0_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_0_V_read[66]);
wire tmp_0_67;
assign tmp_0_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_0_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_0_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_0_V_read[67]);
wire tmp_0_68;
assign tmp_0_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_0_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_0_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_0_V_read[68]);
wire tmp_0_69;
assign tmp_0_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_0_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_0_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_0_V_read[69]);
wire tmp_0_70;
assign tmp_0_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_0_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_0_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_0_V_read[70]);
wire tmp_0_71;
assign tmp_0_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_0_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_0_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_0_V_read[71]);
assign ap_return_0 = {1'b0,tmp_0_1,tmp_0_2,tmp_0_3,tmp_0_4,tmp_0_5,tmp_0_6,1'b0,tmp_0_8,1'b0,tmp_0_10,tmp_0_11,tmp_0_12,tmp_0_13,tmp_0_14,tmp_0_15,tmp_0_16,tmp_0_17,tmp_0_18,tmp_0_19,tmp_0_20,tmp_0_21,tmp_0_22,tmp_0_23,tmp_0_24,tmp_0_25,1'b0,tmp_0_27,tmp_0_28,1'b0,tmp_0_30,1'b0,tmp_0_32,tmp_0_33,tmp_0_34,tmp_0_35,tmp_0_36,tmp_0_37,1'b0,1'b0,tmp_0_40,tmp_0_41,tmp_0_42,tmp_0_43,tmp_0_44,tmp_0_45,tmp_0_46,1'b0,tmp_0_48,tmp_0_49,tmp_0_50,tmp_0_51,tmp_0_52,tmp_0_53,tmp_0_54,tmp_0_55,tmp_0_56,tmp_0_57,tmp_0_58,tmp_0_59,tmp_0_60,tmp_0_61,tmp_0_62,tmp_0_63,tmp_0_64,tmp_0_65,tmp_0_66,tmp_0_67,tmp_0_68,tmp_0_69,tmp_0_70,tmp_0_71};
wire tmp_1_0;
assign tmp_1_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_1_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_1_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_1_V_read[0]);
wire tmp_1_1;
assign tmp_1_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_1_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_1_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_1_V_read[1]);
wire tmp_1_2;
assign tmp_1_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_1_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_1_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_1_V_read[2]);
wire tmp_1_3;
assign tmp_1_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_1_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_1_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_1_V_read[3]);
wire tmp_1_4;
assign tmp_1_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_1_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_1_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_1_V_read[4]);
wire tmp_1_5;
assign tmp_1_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_1_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_1_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_1_V_read[5]);
wire tmp_1_6;
assign tmp_1_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_1_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_1_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_1_V_read[6]);
wire tmp_1_7;
assign tmp_1_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_1_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_1_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_1_V_read[7]);
wire tmp_1_8;
assign tmp_1_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_1_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_1_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_1_V_read[8]);
wire tmp_1_9;
assign tmp_1_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_1_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_1_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_1_V_read[9]);
wire tmp_1_11;
assign tmp_1_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_1_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_1_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_1_V_read[11]);
wire tmp_1_12;
assign tmp_1_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_1_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_1_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_1_V_read[12]);
wire tmp_1_13;
assign tmp_1_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_1_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_1_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_1_V_read[13]);
wire tmp_1_14;
assign tmp_1_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_1_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_1_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_1_V_read[14]);
wire tmp_1_16;
assign tmp_1_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_1_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_1_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_1_V_read[16]);
wire tmp_1_17;
assign tmp_1_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_1_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_1_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_1_V_read[17]);
wire tmp_1_18;
assign tmp_1_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_1_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_1_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_1_V_read[18]);
wire tmp_1_19;
assign tmp_1_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_1_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_1_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_1_V_read[19]);
wire tmp_1_20;
assign tmp_1_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_1_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_1_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_1_V_read[20]);
wire tmp_1_21;
assign tmp_1_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_1_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_1_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_1_V_read[21]);
wire tmp_1_22;
assign tmp_1_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_1_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_1_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_1_V_read[22]);
wire tmp_1_24;
assign tmp_1_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_1_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_1_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_1_V_read[24]);
wire tmp_1_25;
assign tmp_1_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_1_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_1_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_1_V_read[25]);
wire tmp_1_26;
assign tmp_1_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_1_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_1_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_1_V_read[26]);
wire tmp_1_27;
assign tmp_1_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_1_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_1_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_1_V_read[27]);
wire tmp_1_28;
assign tmp_1_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_1_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_1_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_1_V_read[28]);
wire tmp_1_29;
assign tmp_1_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_1_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_1_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_1_V_read[29]);
wire tmp_1_30;
assign tmp_1_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_1_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_1_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_1_V_read[30]);
wire tmp_1_31;
assign tmp_1_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_1_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_1_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_1_V_read[31]);
wire tmp_1_32;
assign tmp_1_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_1_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_1_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_1_V_read[32]);
wire tmp_1_35;
assign tmp_1_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_1_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_1_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_1_V_read[35]);
wire tmp_1_36;
assign tmp_1_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_1_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_1_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_1_V_read[36]);
wire tmp_1_37;
assign tmp_1_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_1_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_1_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_1_V_read[37]);
wire tmp_1_38;
assign tmp_1_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_1_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_1_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_1_V_read[38]);
wire tmp_1_40;
assign tmp_1_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_1_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_1_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_1_V_read[40]);
wire tmp_1_41;
assign tmp_1_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_1_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_1_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_1_V_read[41]);
wire tmp_1_42;
assign tmp_1_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_1_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_1_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_1_V_read[42]);
wire tmp_1_43;
assign tmp_1_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_1_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_1_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_1_V_read[43]);
wire tmp_1_44;
assign tmp_1_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_1_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_1_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_1_V_read[44]);
wire tmp_1_45;
assign tmp_1_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_1_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_1_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_1_V_read[45]);
wire tmp_1_46;
assign tmp_1_46 = (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_1_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_1_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_1_V_read[46]);
wire tmp_1_47;
assign tmp_1_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_1_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_1_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_1_V_read[47]);
wire tmp_1_48;
assign tmp_1_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_1_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_1_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_1_V_read[48]);
wire tmp_1_49;
assign tmp_1_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_1_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_1_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_1_V_read[49]);
wire tmp_1_50;
assign tmp_1_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_1_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_1_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_1_V_read[50]);
wire tmp_1_51;
assign tmp_1_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_1_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_1_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_1_V_read[51]);
wire tmp_1_52;
assign tmp_1_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_1_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_1_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_1_V_read[52]);
wire tmp_1_53;
assign tmp_1_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_1_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_1_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_1_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_1_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_1_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_1_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_1_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_1_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_1_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_1_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_1_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_1_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_1_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_1_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_1_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_1_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_1_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_1_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_1_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_1_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_1_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_1_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_1_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_1_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_1_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_1_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_1_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_1_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_1_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_1_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_1_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_1_V_read[53]);
wire tmp_1_54;
assign tmp_1_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_1_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_1_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_1_V_read[54]);
wire tmp_1_56;
assign tmp_1_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_1_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_1_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_1_V_read[56]);
wire tmp_1_57;
assign tmp_1_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_1_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_1_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_1_V_read[57]);
wire tmp_1_58;
assign tmp_1_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_1_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_1_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_1_V_read[58]);
wire tmp_1_59;
assign tmp_1_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_1_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_1_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_1_V_read[59]);
wire tmp_1_60;
assign tmp_1_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_1_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_1_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_1_V_read[60]);
wire tmp_1_61;
assign tmp_1_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_1_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_1_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_1_V_read[61]);
wire tmp_1_62;
assign tmp_1_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_1_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_1_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_1_V_read[62]);
wire tmp_1_63;
assign tmp_1_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_1_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_1_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_1_V_read[63]);
wire tmp_1_64;
assign tmp_1_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_1_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_1_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_1_V_read[64]);
wire tmp_1_65;
assign tmp_1_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_1_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_1_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_1_V_read[65]);
wire tmp_1_66;
assign tmp_1_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_1_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_1_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_1_V_read[66]);
wire tmp_1_67;
assign tmp_1_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_1_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_1_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_1_V_read[67]);
wire tmp_1_68;
assign tmp_1_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_1_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_1_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_1_V_read[68]);
wire tmp_1_69;
assign tmp_1_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_1_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_1_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_1_V_read[69]);
wire tmp_1_70;
assign tmp_1_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_1_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_1_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_1_V_read[70]);
wire tmp_1_71;
assign tmp_1_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_1_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_1_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_1_V_read[71]);
assign ap_return_1 = {tmp_1_0,tmp_1_1,tmp_1_2,tmp_1_3,tmp_1_4,tmp_1_5,tmp_1_6,tmp_1_7,tmp_1_8,tmp_1_9,1'b0,tmp_1_11,tmp_1_12,tmp_1_13,tmp_1_14,1'b0,tmp_1_16,tmp_1_17,tmp_1_18,tmp_1_19,tmp_1_20,tmp_1_21,tmp_1_22,1'b0,tmp_1_24,tmp_1_25,tmp_1_26,tmp_1_27,tmp_1_28,tmp_1_29,tmp_1_30,tmp_1_31,tmp_1_32,1'b0,1'b0,tmp_1_35,tmp_1_36,tmp_1_37,tmp_1_38,1'b0,tmp_1_40,tmp_1_41,tmp_1_42,tmp_1_43,tmp_1_44,tmp_1_45,tmp_1_46,tmp_1_47,tmp_1_48,tmp_1_49,tmp_1_50,tmp_1_51,tmp_1_52,tmp_1_53,tmp_1_54,1'b0,tmp_1_56,tmp_1_57,tmp_1_58,tmp_1_59,tmp_1_60,tmp_1_61,tmp_1_62,tmp_1_63,tmp_1_64,tmp_1_65,tmp_1_66,tmp_1_67,tmp_1_68,tmp_1_69,tmp_1_70,tmp_1_71};
wire tmp_2_0;
assign tmp_2_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_2_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_2_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_2_V_read[0]);
wire tmp_2_1;
assign tmp_2_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_2_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_2_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_2_V_read[1]);
wire tmp_2_2;
assign tmp_2_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_2_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_2_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_2_V_read[2]);
wire tmp_2_3;
assign tmp_2_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_2_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_2_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_2_V_read[3]);
wire tmp_2_4;
assign tmp_2_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_2_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_2_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_2_V_read[4]);
wire tmp_2_5;
assign tmp_2_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_2_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_2_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_2_V_read[5]);
wire tmp_2_6;
assign tmp_2_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_2_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_2_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_2_V_read[6]);
wire tmp_2_7;
assign tmp_2_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_2_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_2_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_2_V_read[7]);
wire tmp_2_8;
assign tmp_2_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_2_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_2_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_2_V_read[8]);
wire tmp_2_9;
assign tmp_2_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_2_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_2_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_2_V_read[9]);
wire tmp_2_10;
assign tmp_2_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_2_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_2_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_2_V_read[10]);
wire tmp_2_11;
assign tmp_2_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_2_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_2_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_2_V_read[11]);
wire tmp_2_12;
assign tmp_2_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_2_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_2_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_2_V_read[12]);
wire tmp_2_13;
assign tmp_2_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_2_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_2_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_2_V_read[13]);
wire tmp_2_16;
assign tmp_2_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_2_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_2_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_2_V_read[16]);
wire tmp_2_17;
assign tmp_2_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_2_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_2_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_2_V_read[17]);
wire tmp_2_18;
assign tmp_2_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_2_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_2_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_2_V_read[18]);
wire tmp_2_19;
assign tmp_2_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_2_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_2_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_2_V_read[19]);
wire tmp_2_20;
assign tmp_2_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_2_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_2_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_2_V_read[20]);
wire tmp_2_21;
assign tmp_2_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_2_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_2_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_2_V_read[21]);
wire tmp_2_22;
assign tmp_2_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_2_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_2_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_2_V_read[22]);
wire tmp_2_23;
assign tmp_2_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_2_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_2_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_2_V_read[23]);
wire tmp_2_24;
assign tmp_2_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_2_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_2_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_2_V_read[24]);
wire tmp_2_25;
assign tmp_2_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_2_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_2_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_2_V_read[25]);
wire tmp_2_26;
assign tmp_2_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_2_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_2_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_2_V_read[26]);
wire tmp_2_27;
assign tmp_2_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_2_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_2_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_2_V_read[27]);
wire tmp_2_29;
assign tmp_2_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_2_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_2_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_2_V_read[29]);
wire tmp_2_30;
assign tmp_2_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_2_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_2_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_2_V_read[30]);
wire tmp_2_32;
assign tmp_2_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_2_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_2_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_2_V_read[32]);
wire tmp_2_33;
assign tmp_2_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_2_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_2_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_2_V_read[33]);
wire tmp_2_34;
assign tmp_2_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_2_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_2_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_2_V_read[34]);
wire tmp_2_35;
assign tmp_2_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_2_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_2_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_2_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_2_V_read[35]);
wire tmp_2_36;
assign tmp_2_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_2_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_2_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_2_V_read[36]);
wire tmp_2_37;
assign tmp_2_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_2_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_2_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_2_V_read[37]);
wire tmp_2_38;
assign tmp_2_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_2_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_2_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_2_V_read[38]);
wire tmp_2_39;
assign tmp_2_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_2_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_2_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_2_V_read[39]);
wire tmp_2_40;
assign tmp_2_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_2_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_2_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_2_V_read[40]);
wire tmp_2_41;
assign tmp_2_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_2_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_2_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_2_V_read[41]);
wire tmp_2_42;
assign tmp_2_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_2_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_2_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_2_V_read[42]);
wire tmp_2_43;
assign tmp_2_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_2_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_2_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_2_V_read[43]);
wire tmp_2_44;
assign tmp_2_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_2_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_2_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_2_V_read[44]);
wire tmp_2_45;
assign tmp_2_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_2_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_2_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_2_V_read[45]);
wire tmp_2_46;
assign tmp_2_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_2_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_2_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_2_V_read[46]);
wire tmp_2_48;
assign tmp_2_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_2_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_2_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_2_V_read[48]);
wire tmp_2_49;
assign tmp_2_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_2_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_2_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_2_V_read[49]);
wire tmp_2_50;
assign tmp_2_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_2_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_2_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_2_V_read[50]);
wire tmp_2_51;
assign tmp_2_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_2_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_2_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_2_V_read[51]);
wire tmp_2_52;
assign tmp_2_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_2_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_2_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_2_V_read[52]);
wire tmp_2_54;
assign tmp_2_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_2_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_2_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_2_V_read[54]);
wire tmp_2_56;
assign tmp_2_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_2_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_2_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_2_V_read[56]);
wire tmp_2_57;
assign tmp_2_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_2_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_2_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_2_V_read[57]);
wire tmp_2_59;
assign tmp_2_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_2_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_2_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_2_V_read[59]);
wire tmp_2_60;
assign tmp_2_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_2_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_2_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_2_V_read[60]);
wire tmp_2_61;
assign tmp_2_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_2_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_2_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_2_V_read[61]);
wire tmp_2_62;
assign tmp_2_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_2_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_2_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_2_V_read[62]);
wire tmp_2_63;
assign tmp_2_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_2_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_2_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_2_V_read[63]);
wire tmp_2_66;
assign tmp_2_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_2_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_2_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_2_V_read[66]);
wire tmp_2_67;
assign tmp_2_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_2_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_2_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_2_V_read[67]);
wire tmp_2_68;
assign tmp_2_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_2_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_2_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_2_V_read[68]);
wire tmp_2_69;
assign tmp_2_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_2_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_2_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_2_V_read[69]);
wire tmp_2_70;
assign tmp_2_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_2_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_2_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_2_V_read[70]);
wire tmp_2_71;
assign tmp_2_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_2_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_2_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_2_V_read[71]);
assign ap_return_2 = {tmp_2_0,tmp_2_1,tmp_2_2,tmp_2_3,tmp_2_4,tmp_2_5,tmp_2_6,tmp_2_7,tmp_2_8,tmp_2_9,tmp_2_10,tmp_2_11,tmp_2_12,tmp_2_13,1'b0,1'b0,tmp_2_16,tmp_2_17,tmp_2_18,tmp_2_19,tmp_2_20,tmp_2_21,tmp_2_22,tmp_2_23,tmp_2_24,tmp_2_25,tmp_2_26,tmp_2_27,1'b0,tmp_2_29,tmp_2_30,1'b0,tmp_2_32,tmp_2_33,tmp_2_34,tmp_2_35,tmp_2_36,tmp_2_37,tmp_2_38,tmp_2_39,tmp_2_40,tmp_2_41,tmp_2_42,tmp_2_43,tmp_2_44,tmp_2_45,tmp_2_46,1'b0,tmp_2_48,tmp_2_49,tmp_2_50,tmp_2_51,tmp_2_52,1'b0,tmp_2_54,1'b0,tmp_2_56,tmp_2_57,1'b0,tmp_2_59,tmp_2_60,tmp_2_61,tmp_2_62,tmp_2_63,1'b0,1'b0,tmp_2_66,tmp_2_67,tmp_2_68,tmp_2_69,tmp_2_70,tmp_2_71};
wire tmp_3_0;
assign tmp_3_0 = (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_3_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_3_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_3_V_read[0]);
wire tmp_3_1;
assign tmp_3_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_3_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_3_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_3_V_read[1]);
wire tmp_3_2;
assign tmp_3_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_3_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_3_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_3_V_read[2]);
wire tmp_3_3;
assign tmp_3_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_3_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_3_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_3_V_read[3]);
wire tmp_3_4;
assign tmp_3_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_3_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_3_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_3_V_read[4]);
wire tmp_3_5;
assign tmp_3_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_3_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_3_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_3_V_read[5]);
wire tmp_3_6;
assign tmp_3_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_3_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_3_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_3_V_read[6]);
wire tmp_3_7;
assign tmp_3_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_3_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_3_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_3_V_read[7]);
wire tmp_3_8;
assign tmp_3_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_3_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_3_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_3_V_read[8]);
wire tmp_3_9;
assign tmp_3_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_3_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_3_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_3_V_read[9]);
wire tmp_3_11;
assign tmp_3_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_3_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_3_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_3_V_read[11]);
wire tmp_3_12;
assign tmp_3_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_3_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_3_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_3_V_read[12]);
wire tmp_3_13;
assign tmp_3_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_3_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_3_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_3_V_read[13]);
wire tmp_3_14;
assign tmp_3_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_3_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_3_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_3_V_read[14]);
wire tmp_3_16;
assign tmp_3_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_3_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_3_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_3_V_read[16]);
wire tmp_3_17;
assign tmp_3_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_3_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_3_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_3_V_read[17]);
wire tmp_3_18;
assign tmp_3_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_3_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_3_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_3_V_read[18]);
wire tmp_3_19;
assign tmp_3_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_3_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_3_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_3_V_read[19]);
wire tmp_3_20;
assign tmp_3_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_3_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_3_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_3_V_read[20]);
wire tmp_3_21;
assign tmp_3_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_3_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_3_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_3_V_read[21]);
wire tmp_3_22;
assign tmp_3_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_3_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_3_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_3_V_read[22]);
wire tmp_3_23;
assign tmp_3_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_3_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_3_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_3_V_read[23]);
wire tmp_3_24;
assign tmp_3_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_3_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_3_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_3_V_read[24]);
wire tmp_3_25;
assign tmp_3_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_3_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_3_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_3_V_read[25]);
wire tmp_3_26;
assign tmp_3_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_3_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_3_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_3_V_read[26]);
wire tmp_3_27;
assign tmp_3_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_3_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_3_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_3_V_read[27]);
wire tmp_3_28;
assign tmp_3_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_3_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_3_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_3_V_read[28]);
wire tmp_3_29;
assign tmp_3_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_3_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_3_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_3_V_read[29]);
wire tmp_3_30;
assign tmp_3_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_3_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_3_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_3_V_read[30]);
wire tmp_3_32;
assign tmp_3_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_3_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_3_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_3_V_read[32]);
wire tmp_3_33;
assign tmp_3_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_3_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_3_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_3_V_read[33]);
wire tmp_3_35;
assign tmp_3_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_3_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_3_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_3_V_read[35]);
wire tmp_3_36;
assign tmp_3_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_3_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_3_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_3_V_read[36]);
wire tmp_3_38;
assign tmp_3_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_3_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_3_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_3_V_read[38]);
wire tmp_3_40;
assign tmp_3_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_3_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_3_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_3_V_read[40]);
wire tmp_3_41;
assign tmp_3_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_3_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_3_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_3_V_read[41]);
wire tmp_3_42;
assign tmp_3_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_3_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_3_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_3_V_read[42]);
wire tmp_3_45;
assign tmp_3_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_3_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_3_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_3_V_read[45]);
wire tmp_3_49;
assign tmp_3_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_3_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_3_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_3_V_read[49]);
wire tmp_3_50;
assign tmp_3_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_3_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_3_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_3_V_read[50]);
wire tmp_3_51;
assign tmp_3_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_3_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_3_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_3_V_read[51]);
wire tmp_3_52;
assign tmp_3_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_3_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_3_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_3_V_read[52]);
wire tmp_3_53;
assign tmp_3_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_3_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_3_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_3_V_read[53]);
wire tmp_3_54;
assign tmp_3_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_3_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_3_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_3_V_read[54]);
wire tmp_3_55;
assign tmp_3_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_3_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_3_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_3_V_read[55]);
wire tmp_3_56;
assign tmp_3_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_3_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_3_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_3_V_read[56]);
wire tmp_3_57;
assign tmp_3_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_3_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_3_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_3_V_read[57]);
wire tmp_3_59;
assign tmp_3_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_3_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_3_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_3_V_read[59]);
wire tmp_3_61;
assign tmp_3_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_3_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_3_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_3_V_read[61]);
wire tmp_3_62;
assign tmp_3_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_3_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_3_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_3_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_3_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_3_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_3_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_3_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_3_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_3_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_3_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_3_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_3_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_3_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_3_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_3_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_3_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_3_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_3_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_3_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_3_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_3_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_3_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_3_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_3_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_3_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_3_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_3_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_3_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_3_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_3_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_3_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_3_V_read[62]);
wire tmp_3_63;
assign tmp_3_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_3_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_3_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_3_V_read[63]);
wire tmp_3_65;
assign tmp_3_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_3_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_3_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_3_V_read[65]);
wire tmp_3_66;
assign tmp_3_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_3_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_3_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_3_V_read[66]);
wire tmp_3_67;
assign tmp_3_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_3_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_3_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_3_V_read[67]);
wire tmp_3_68;
assign tmp_3_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_3_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_3_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_3_V_read[68]);
wire tmp_3_70;
assign tmp_3_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_3_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_3_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_3_V_read[70]);
wire tmp_3_71;
assign tmp_3_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_3_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_3_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_3_V_read[71]);
assign ap_return_3 = {tmp_3_0,tmp_3_1,tmp_3_2,tmp_3_3,tmp_3_4,tmp_3_5,tmp_3_6,tmp_3_7,tmp_3_8,tmp_3_9,1'b0,tmp_3_11,tmp_3_12,tmp_3_13,tmp_3_14,1'b0,tmp_3_16,tmp_3_17,tmp_3_18,tmp_3_19,tmp_3_20,tmp_3_21,tmp_3_22,tmp_3_23,tmp_3_24,tmp_3_25,tmp_3_26,tmp_3_27,tmp_3_28,tmp_3_29,tmp_3_30,1'b0,tmp_3_32,tmp_3_33,1'b0,tmp_3_35,tmp_3_36,1'b0,tmp_3_38,1'b0,tmp_3_40,tmp_3_41,tmp_3_42,1'b0,1'b0,tmp_3_45,1'b0,1'b0,1'b0,tmp_3_49,tmp_3_50,tmp_3_51,tmp_3_52,tmp_3_53,tmp_3_54,tmp_3_55,tmp_3_56,tmp_3_57,1'b0,tmp_3_59,1'b0,tmp_3_61,tmp_3_62,tmp_3_63,1'b0,tmp_3_65,tmp_3_66,tmp_3_67,tmp_3_68,1'b0,tmp_3_70,tmp_3_71};
wire tmp_4_0;
assign tmp_4_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_4_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_4_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_4_V_read[0]);
wire tmp_4_1;
assign tmp_4_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_4_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_4_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_4_V_read[1]);
wire tmp_4_2;
assign tmp_4_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_4_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_4_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_4_V_read[2]);
wire tmp_4_3;
assign tmp_4_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_4_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_4_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_4_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_4_V_read[3]);
wire tmp_4_4;
assign tmp_4_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_4_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_4_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_4_V_read[4]);
wire tmp_4_5;
assign tmp_4_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_4_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_4_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_4_V_read[5]);
wire tmp_4_6;
assign tmp_4_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_4_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_4_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_4_V_read[6]);
wire tmp_4_7;
assign tmp_4_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_4_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_4_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_4_V_read[7]);
wire tmp_4_8;
assign tmp_4_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_4_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_4_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_4_V_read[8]);
wire tmp_4_9;
assign tmp_4_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_4_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_4_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_4_V_read[9]);
wire tmp_4_11;
assign tmp_4_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_4_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_4_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_4_V_read[11]);
wire tmp_4_12;
assign tmp_4_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_4_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_4_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_4_V_read[12]);
wire tmp_4_13;
assign tmp_4_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_4_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_4_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_4_V_read[13]);
wire tmp_4_14;
assign tmp_4_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_4_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_4_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_4_V_read[14]);
wire tmp_4_16;
assign tmp_4_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_4_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_4_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_4_V_read[16]);
wire tmp_4_17;
assign tmp_4_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_4_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_4_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_4_V_read[17]);
wire tmp_4_18;
assign tmp_4_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_4_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_4_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_4_V_read[18]);
wire tmp_4_19;
assign tmp_4_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_4_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_4_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_4_V_read[19]);
wire tmp_4_20;
assign tmp_4_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_4_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_4_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_4_V_read[20]);
wire tmp_4_21;
assign tmp_4_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_4_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_4_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_4_V_read[21]);
wire tmp_4_22;
assign tmp_4_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_4_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_4_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_4_V_read[22]);
wire tmp_4_23;
assign tmp_4_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_4_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_4_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_4_V_read[23]);
wire tmp_4_24;
assign tmp_4_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_4_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_4_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_4_V_read[24]);
wire tmp_4_26;
assign tmp_4_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_4_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_4_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_4_V_read[26]);
wire tmp_4_27;
assign tmp_4_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_4_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_4_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_4_V_read[27]);
wire tmp_4_28;
assign tmp_4_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_4_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_4_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_4_V_read[28]);
wire tmp_4_29;
assign tmp_4_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_4_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_4_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_4_V_read[29]);
wire tmp_4_30;
assign tmp_4_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_4_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_4_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_4_V_read[30]);
wire tmp_4_31;
assign tmp_4_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_4_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_4_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_4_V_read[31]);
wire tmp_4_32;
assign tmp_4_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_4_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_4_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_4_V_read[32]);
wire tmp_4_33;
assign tmp_4_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_4_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_4_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_4_V_read[33]);
wire tmp_4_34;
assign tmp_4_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_4_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_4_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_4_V_read[34]);
wire tmp_4_35;
assign tmp_4_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_4_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_4_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_4_V_read[35]);
wire tmp_4_36;
assign tmp_4_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_4_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_4_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_4_V_read[36]);
wire tmp_4_37;
assign tmp_4_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_4_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_4_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_4_V_read[37]);
wire tmp_4_38;
assign tmp_4_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_4_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_4_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_4_V_read[38]);
wire tmp_4_39;
assign tmp_4_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_4_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_4_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_4_V_read[39]);
wire tmp_4_40;
assign tmp_4_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_4_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_4_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_4_V_read[40]);
wire tmp_4_41;
assign tmp_4_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_4_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_4_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_4_V_read[41]);
wire tmp_4_42;
assign tmp_4_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_4_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_4_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_4_V_read[42]);
wire tmp_4_43;
assign tmp_4_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_4_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_4_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_4_V_read[43]);
wire tmp_4_44;
assign tmp_4_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_4_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_4_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_4_V_read[44]);
wire tmp_4_45;
assign tmp_4_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_4_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_4_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_4_V_read[45]);
wire tmp_4_47;
assign tmp_4_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_4_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_4_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_4_V_read[47]);
wire tmp_4_48;
assign tmp_4_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_4_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_4_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_4_V_read[48]);
wire tmp_4_49;
assign tmp_4_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_4_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_4_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_4_V_read[49]);
wire tmp_4_50;
assign tmp_4_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_4_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_4_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_4_V_read[50]);
wire tmp_4_51;
assign tmp_4_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_4_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_4_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_4_V_read[51]);
wire tmp_4_52;
assign tmp_4_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_4_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_4_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_4_V_read[52]);
wire tmp_4_53;
assign tmp_4_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_4_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_4_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_4_V_read[53]);
wire tmp_4_54;
assign tmp_4_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_4_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_4_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_4_V_read[54]);
wire tmp_4_55;
assign tmp_4_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_4_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_4_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_4_V_read[55]);
wire tmp_4_56;
assign tmp_4_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_4_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_4_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_4_V_read[56]);
wire tmp_4_57;
assign tmp_4_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_4_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_4_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_4_V_read[57]);
wire tmp_4_58;
assign tmp_4_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_4_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_4_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_4_V_read[58]);
wire tmp_4_59;
assign tmp_4_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_4_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_4_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_4_V_read[59]);
wire tmp_4_60;
assign tmp_4_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_4_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_4_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_4_V_read[60]);
wire tmp_4_61;
assign tmp_4_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_4_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_4_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_4_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_4_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_4_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_4_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_4_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_4_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_4_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_4_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_4_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_4_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_4_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_4_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_4_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_4_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_4_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_4_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_4_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_4_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_4_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_4_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_4_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_4_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_4_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_4_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_4_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_4_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_4_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_4_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_4_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_4_V_read[61]);
wire tmp_4_63;
assign tmp_4_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_4_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_4_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_4_V_read[63]);
wire tmp_4_64;
assign tmp_4_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_4_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_4_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_4_V_read[64]);
wire tmp_4_65;
assign tmp_4_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_4_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_4_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_4_V_read[65]);
wire tmp_4_66;
assign tmp_4_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_4_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_4_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_4_V_read[66]);
wire tmp_4_67;
assign tmp_4_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_4_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_4_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_4_V_read[67]);
wire tmp_4_68;
assign tmp_4_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_4_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_4_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_4_V_read[68]);
wire tmp_4_69;
assign tmp_4_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_4_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_4_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_4_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_4_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_4_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_4_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_4_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_4_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_4_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_4_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_4_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_4_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_4_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_4_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_4_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_4_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_4_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_4_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_4_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_4_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_4_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_4_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_4_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_4_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_4_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_4_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_4_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_4_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_4_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_4_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_4_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_4_V_read[69]);
wire tmp_4_70;
assign tmp_4_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_4_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_4_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_4_V_read[70]);
assign ap_return_4 = {tmp_4_0,tmp_4_1,tmp_4_2,tmp_4_3,tmp_4_4,tmp_4_5,tmp_4_6,tmp_4_7,tmp_4_8,tmp_4_9,1'b0,tmp_4_11,tmp_4_12,tmp_4_13,tmp_4_14,1'b0,tmp_4_16,tmp_4_17,tmp_4_18,tmp_4_19,tmp_4_20,tmp_4_21,tmp_4_22,tmp_4_23,tmp_4_24,1'b0,tmp_4_26,tmp_4_27,tmp_4_28,tmp_4_29,tmp_4_30,tmp_4_31,tmp_4_32,tmp_4_33,tmp_4_34,tmp_4_35,tmp_4_36,tmp_4_37,tmp_4_38,tmp_4_39,tmp_4_40,tmp_4_41,tmp_4_42,tmp_4_43,tmp_4_44,tmp_4_45,1'b0,tmp_4_47,tmp_4_48,tmp_4_49,tmp_4_50,tmp_4_51,tmp_4_52,tmp_4_53,tmp_4_54,tmp_4_55,tmp_4_56,tmp_4_57,tmp_4_58,tmp_4_59,tmp_4_60,tmp_4_61,1'b0,tmp_4_63,tmp_4_64,tmp_4_65,tmp_4_66,tmp_4_67,tmp_4_68,tmp_4_69,tmp_4_70,1'b0};
wire tmp_5_0;
assign tmp_5_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_5_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_5_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_5_V_read[0]);
wire tmp_5_1;
assign tmp_5_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_5_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_5_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_5_V_read[1]);
wire tmp_5_2;
assign tmp_5_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_5_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_5_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_5_V_read[2]);
wire tmp_5_3;
assign tmp_5_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_5_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_5_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_5_V_read[3]);
wire tmp_5_4;
assign tmp_5_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_5_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_5_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_5_V_read[4]);
wire tmp_5_5;
assign tmp_5_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_5_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_5_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_5_V_read[5]);
wire tmp_5_6;
assign tmp_5_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_5_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_5_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_5_V_read[6]);
wire tmp_5_7;
assign tmp_5_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_5_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_5_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_5_V_read[7]);
wire tmp_5_8;
assign tmp_5_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_5_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_5_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_5_V_read[8]);
wire tmp_5_9;
assign tmp_5_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_5_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_5_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_5_V_read[9]);
wire tmp_5_10;
assign tmp_5_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_5_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_5_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_5_V_read[10]);
wire tmp_5_11;
assign tmp_5_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_5_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_5_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_5_V_read[11]);
wire tmp_5_12;
assign tmp_5_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_5_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_5_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_5_V_read[12]);
wire tmp_5_13;
assign tmp_5_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_5_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_5_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_5_V_read[13]);
wire tmp_5_16;
assign tmp_5_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_5_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_5_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_5_V_read[16]);
wire tmp_5_17;
assign tmp_5_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_5_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_5_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_5_V_read[17]);
wire tmp_5_18;
assign tmp_5_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_5_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_5_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_5_V_read[18]);
wire tmp_5_19;
assign tmp_5_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_5_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_5_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_5_V_read[19]);
wire tmp_5_20;
assign tmp_5_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_5_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_5_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_5_V_read[20]);
wire tmp_5_21;
assign tmp_5_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_5_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_5_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_5_V_read[21]);
wire tmp_5_22;
assign tmp_5_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_5_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_5_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_5_V_read[22]);
wire tmp_5_23;
assign tmp_5_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_5_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_5_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_5_V_read[23]);
wire tmp_5_24;
assign tmp_5_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_5_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_5_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_5_V_read[24]);
wire tmp_5_25;
assign tmp_5_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_5_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_5_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_5_V_read[25]);
wire tmp_5_26;
assign tmp_5_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_5_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_5_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_5_V_read[26]);
wire tmp_5_27;
assign tmp_5_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_5_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_5_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_5_V_read[27]);
wire tmp_5_28;
assign tmp_5_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_5_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_5_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_5_V_read[28]);
wire tmp_5_29;
assign tmp_5_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_5_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_5_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_5_V_read[29]);
wire tmp_5_30;
assign tmp_5_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_5_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_5_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_5_V_read[30]);
wire tmp_5_31;
assign tmp_5_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_5_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_5_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_5_V_read[31]);
wire tmp_5_32;
assign tmp_5_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_5_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_5_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_5_V_read[32]);
wire tmp_5_33;
assign tmp_5_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_5_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_5_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_5_V_read[33]);
wire tmp_5_35;
assign tmp_5_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_5_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_5_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_5_V_read[35]);
wire tmp_5_36;
assign tmp_5_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_5_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_5_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_5_V_read[36]);
wire tmp_5_37;
assign tmp_5_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_5_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_5_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_5_V_read[37]);
wire tmp_5_38;
assign tmp_5_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_5_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_5_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_5_V_read[38]);
wire tmp_5_40;
assign tmp_5_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_5_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_5_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_5_V_read[40]);
wire tmp_5_41;
assign tmp_5_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_5_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_5_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_5_V_read[41]);
wire tmp_5_42;
assign tmp_5_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_5_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_5_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_5_V_read[42]);
wire tmp_5_43;
assign tmp_5_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_5_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_5_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_5_V_read[43]);
wire tmp_5_44;
assign tmp_5_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_5_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_5_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_5_V_read[44]);
wire tmp_5_45;
assign tmp_5_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_5_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_5_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_5_V_read[45]);
wire tmp_5_47;
assign tmp_5_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_5_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_5_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_5_V_read[47]);
wire tmp_5_48;
assign tmp_5_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_5_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_5_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_5_V_read[48]);
wire tmp_5_49;
assign tmp_5_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_5_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_5_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_5_V_read[49]);
wire tmp_5_50;
assign tmp_5_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_5_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_5_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_5_V_read[50]);
wire tmp_5_51;
assign tmp_5_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_5_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_5_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_5_V_read[51]);
wire tmp_5_52;
assign tmp_5_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_5_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_5_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_5_V_read[52]);
wire tmp_5_53;
assign tmp_5_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_5_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_5_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_5_V_read[53]);
wire tmp_5_54;
assign tmp_5_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_5_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_5_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_5_V_read[54]);
wire tmp_5_55;
assign tmp_5_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_5_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_5_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_5_V_read[55]);
wire tmp_5_56;
assign tmp_5_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_5_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_5_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_5_V_read[56]);
wire tmp_5_57;
assign tmp_5_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_5_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_5_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_5_V_read[57]);
wire tmp_5_59;
assign tmp_5_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_5_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_5_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_5_V_read[59]);
wire tmp_5_60;
assign tmp_5_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_5_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_5_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_5_V_read[60]);
wire tmp_5_61;
assign tmp_5_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_5_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_5_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_5_V_read[61]);
wire tmp_5_62;
assign tmp_5_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_5_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_5_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_5_V_read[62]);
wire tmp_5_63;
assign tmp_5_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_5_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_5_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_5_V_read[63]);
wire tmp_5_64;
assign tmp_5_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_5_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_5_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_5_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_5_V_read[64]);
wire tmp_5_65;
assign tmp_5_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_5_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_5_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_5_V_read[65]);
wire tmp_5_66;
assign tmp_5_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_5_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_5_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_5_V_read[66]);
wire tmp_5_67;
assign tmp_5_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_5_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_5_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_5_V_read[67]);
wire tmp_5_68;
assign tmp_5_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_5_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_5_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_5_V_read[68]);
wire tmp_5_69;
assign tmp_5_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_5_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_5_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_5_V_read[69]);
wire tmp_5_70;
assign tmp_5_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_5_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_5_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_5_V_read[70]);
wire tmp_5_71;
assign tmp_5_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_5_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_5_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_5_V_read[71]);
assign ap_return_5 = {tmp_5_0,tmp_5_1,tmp_5_2,tmp_5_3,tmp_5_4,tmp_5_5,tmp_5_6,tmp_5_7,tmp_5_8,tmp_5_9,tmp_5_10,tmp_5_11,tmp_5_12,tmp_5_13,1'b0,1'b0,tmp_5_16,tmp_5_17,tmp_5_18,tmp_5_19,tmp_5_20,tmp_5_21,tmp_5_22,tmp_5_23,tmp_5_24,tmp_5_25,tmp_5_26,tmp_5_27,tmp_5_28,tmp_5_29,tmp_5_30,tmp_5_31,tmp_5_32,tmp_5_33,1'b0,tmp_5_35,tmp_5_36,tmp_5_37,tmp_5_38,1'b0,tmp_5_40,tmp_5_41,tmp_5_42,tmp_5_43,tmp_5_44,tmp_5_45,1'b0,tmp_5_47,tmp_5_48,tmp_5_49,tmp_5_50,tmp_5_51,tmp_5_52,tmp_5_53,tmp_5_54,tmp_5_55,tmp_5_56,tmp_5_57,1'b0,tmp_5_59,tmp_5_60,tmp_5_61,tmp_5_62,tmp_5_63,tmp_5_64,tmp_5_65,tmp_5_66,tmp_5_67,tmp_5_68,tmp_5_69,tmp_5_70,tmp_5_71};
wire tmp_6_0;
assign tmp_6_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_6_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_6_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_6_V_read[0]);
wire tmp_6_1;
assign tmp_6_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_6_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_6_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_6_V_read[1]);
wire tmp_6_2;
assign tmp_6_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_6_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_6_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_6_V_read[2]);
wire tmp_6_3;
assign tmp_6_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_6_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_6_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_6_V_read[3]);
wire tmp_6_4;
assign tmp_6_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_6_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_6_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_6_V_read[4]);
wire tmp_6_5;
assign tmp_6_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_6_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_6_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_6_V_read[5]);
wire tmp_6_6;
assign tmp_6_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_6_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_6_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_6_V_read[6]);
wire tmp_6_9;
assign tmp_6_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_6_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_6_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_6_V_read[9]);
wire tmp_6_10;
assign tmp_6_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_6_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_6_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_6_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_6_V_read[10]);
wire tmp_6_11;
assign tmp_6_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_6_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_6_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_6_V_read[11]);
wire tmp_6_12;
assign tmp_6_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_6_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_6_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_6_V_read[12]);
wire tmp_6_13;
assign tmp_6_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_6_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_6_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_6_V_read[13]);
wire tmp_6_14;
assign tmp_6_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_6_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_6_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_6_V_read[14]);
wire tmp_6_15;
assign tmp_6_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_6_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_6_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_6_V_read[15]);
wire tmp_6_16;
assign tmp_6_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_6_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_6_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_6_V_read[16]);
wire tmp_6_17;
assign tmp_6_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_6_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_6_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_6_V_read[17]);
wire tmp_6_18;
assign tmp_6_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_6_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_6_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_6_V_read[18]);
wire tmp_6_19;
assign tmp_6_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_6_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_6_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_6_V_read[19]);
wire tmp_6_20;
assign tmp_6_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_6_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_6_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_6_V_read[20]);
wire tmp_6_21;
assign tmp_6_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_6_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_6_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_6_V_read[21]);
wire tmp_6_22;
assign tmp_6_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_6_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_6_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_6_V_read[22]);
wire tmp_6_24;
assign tmp_6_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_6_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_6_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_6_V_read[24]);
wire tmp_6_25;
assign tmp_6_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_6_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_6_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_6_V_read[25]);
wire tmp_6_26;
assign tmp_6_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_6_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_6_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_6_V_read[26]);
wire tmp_6_27;
assign tmp_6_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_6_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_6_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_6_V_read[27]);
wire tmp_6_28;
assign tmp_6_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_6_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_6_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_6_V_read[28]);
wire tmp_6_29;
assign tmp_6_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_6_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_6_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_6_V_read[29]);
wire tmp_6_30;
assign tmp_6_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_6_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_6_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_6_V_read[30]);
wire tmp_6_31;
assign tmp_6_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_6_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_6_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_6_V_read[31]);
wire tmp_6_32;
assign tmp_6_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_6_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_6_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_6_V_read[32]);
wire tmp_6_33;
assign tmp_6_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_6_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_6_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_6_V_read[33]);
wire tmp_6_36;
assign tmp_6_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_6_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_6_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_6_V_read[36]);
wire tmp_6_37;
assign tmp_6_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_6_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_6_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_6_V_read[37]);
wire tmp_6_38;
assign tmp_6_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_6_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_6_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_6_V_read[38]);
wire tmp_6_39;
assign tmp_6_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_6_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_6_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_6_V_read[39]);
wire tmp_6_40;
assign tmp_6_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_6_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_6_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_6_V_read[40]);
wire tmp_6_41;
assign tmp_6_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_6_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_6_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_6_V_read[41]);
wire tmp_6_42;
assign tmp_6_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_6_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_6_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_6_V_read[42]);
wire tmp_6_43;
assign tmp_6_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_6_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_6_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_6_V_read[43]);
wire tmp_6_44;
assign tmp_6_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_6_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_6_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_6_V_read[44]);
wire tmp_6_45;
assign tmp_6_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_6_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_6_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_6_V_read[45]);
wire tmp_6_46;
assign tmp_6_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_6_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_6_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_6_V_read[46]);
wire tmp_6_47;
assign tmp_6_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_6_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_6_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_6_V_read[47]);
wire tmp_6_48;
assign tmp_6_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_6_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_6_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_6_V_read[48]);
wire tmp_6_49;
assign tmp_6_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_6_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_6_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_6_V_read[49]);
wire tmp_6_50;
assign tmp_6_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_6_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_6_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_6_V_read[50]);
wire tmp_6_51;
assign tmp_6_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_6_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_6_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_6_V_read[51]);
wire tmp_6_52;
assign tmp_6_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_6_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_6_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_6_V_read[52]);
wire tmp_6_53;
assign tmp_6_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_6_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_6_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_6_V_read[53]);
wire tmp_6_55;
assign tmp_6_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_6_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_6_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_6_V_read[55]);
wire tmp_6_56;
assign tmp_6_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_6_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_6_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_6_V_read[56]);
wire tmp_6_57;
assign tmp_6_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_6_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_6_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_6_V_read[57]);
wire tmp_6_58;
assign tmp_6_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_6_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_6_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_6_V_read[58]);
wire tmp_6_59;
assign tmp_6_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_6_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_6_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_6_V_read[59]);
wire tmp_6_60;
assign tmp_6_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_6_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_6_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_6_V_read[60]);
wire tmp_6_61;
assign tmp_6_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_6_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_6_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_6_V_read[61]);
wire tmp_6_63;
assign tmp_6_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_6_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_6_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_6_V_read[63]);
wire tmp_6_64;
assign tmp_6_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_6_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_6_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_6_V_read[64]);
wire tmp_6_65;
assign tmp_6_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_6_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_6_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_6_V_read[65]);
wire tmp_6_66;
assign tmp_6_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_6_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_6_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_6_V_read[66]);
wire tmp_6_67;
assign tmp_6_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_6_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_6_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_6_V_read[67]);
wire tmp_6_68;
assign tmp_6_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_6_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_6_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_6_V_read[68]);
wire tmp_6_69;
assign tmp_6_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_6_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_6_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_6_V_read[69]);
wire tmp_6_70;
assign tmp_6_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_6_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_6_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_6_V_read[70]);
wire tmp_6_71;
assign tmp_6_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_6_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_6_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_6_V_read[71]);
assign ap_return_6 = {tmp_6_0,tmp_6_1,tmp_6_2,tmp_6_3,tmp_6_4,tmp_6_5,tmp_6_6,1'b0,1'b0,tmp_6_9,tmp_6_10,tmp_6_11,tmp_6_12,tmp_6_13,tmp_6_14,tmp_6_15,tmp_6_16,tmp_6_17,tmp_6_18,tmp_6_19,tmp_6_20,tmp_6_21,tmp_6_22,1'b0,tmp_6_24,tmp_6_25,tmp_6_26,tmp_6_27,tmp_6_28,tmp_6_29,tmp_6_30,tmp_6_31,tmp_6_32,tmp_6_33,1'b0,1'b0,tmp_6_36,tmp_6_37,tmp_6_38,tmp_6_39,tmp_6_40,tmp_6_41,tmp_6_42,tmp_6_43,tmp_6_44,tmp_6_45,tmp_6_46,tmp_6_47,tmp_6_48,tmp_6_49,tmp_6_50,tmp_6_51,tmp_6_52,tmp_6_53,1'b0,tmp_6_55,tmp_6_56,tmp_6_57,tmp_6_58,tmp_6_59,tmp_6_60,tmp_6_61,1'b0,tmp_6_63,tmp_6_64,tmp_6_65,tmp_6_66,tmp_6_67,tmp_6_68,tmp_6_69,tmp_6_70,tmp_6_71};
wire tmp_7_0;
assign tmp_7_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_7_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_7_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_7_V_read[0]);
wire tmp_7_1;
assign tmp_7_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_7_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_7_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_7_V_read[1]);
wire tmp_7_2;
assign tmp_7_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_7_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_7_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_7_V_read[2]);
wire tmp_7_3;
assign tmp_7_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_7_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_7_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_7_V_read[3]);
wire tmp_7_4;
assign tmp_7_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_7_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_7_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_7_V_read[4]);
wire tmp_7_5;
assign tmp_7_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_7_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_7_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_7_V_read[5]);
wire tmp_7_6;
assign tmp_7_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_7_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_7_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_7_V_read[6]);
wire tmp_7_7;
assign tmp_7_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_7_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_7_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_7_V_read[7]);
wire tmp_7_9;
assign tmp_7_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_7_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_7_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_7_V_read[9]);
wire tmp_7_10;
assign tmp_7_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_7_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_7_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_7_V_read[10]);
wire tmp_7_12;
assign tmp_7_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_7_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_7_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_7_V_read[12]);
wire tmp_7_13;
assign tmp_7_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_7_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_7_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_7_V_read[13]);
wire tmp_7_14;
assign tmp_7_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_7_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_7_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_7_V_read[14]);
wire tmp_7_15;
assign tmp_7_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_7_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_7_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_7_V_read[15]);
wire tmp_7_16;
assign tmp_7_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_7_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_7_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_7_V_read[16]);
wire tmp_7_17;
assign tmp_7_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_7_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_7_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_7_V_read[17]);
wire tmp_7_18;
assign tmp_7_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_7_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_7_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_7_V_read[18]);
wire tmp_7_19;
assign tmp_7_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_7_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_7_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_7_V_read[19]);
wire tmp_7_20;
assign tmp_7_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_7_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_7_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_7_V_read[20]);
wire tmp_7_21;
assign tmp_7_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_7_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_7_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_7_V_read[21]);
wire tmp_7_22;
assign tmp_7_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_7_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_7_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_7_V_read[22]);
wire tmp_7_23;
assign tmp_7_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_7_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_7_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_7_V_read[23]);
wire tmp_7_24;
assign tmp_7_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_7_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_7_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_7_V_read[24]);
wire tmp_7_26;
assign tmp_7_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_7_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_7_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_7_V_read[26]);
wire tmp_7_27;
assign tmp_7_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_7_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_7_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_7_V_read[27]);
wire tmp_7_28;
assign tmp_7_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_7_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_7_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_7_V_read[28]);
wire tmp_7_29;
assign tmp_7_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_7_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_7_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_7_V_read[29]);
wire tmp_7_30;
assign tmp_7_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_7_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_7_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_7_V_read[30]);
wire tmp_7_31;
assign tmp_7_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_7_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_7_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_7_V_read[31]);
wire tmp_7_32;
assign tmp_7_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_7_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_7_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_7_V_read[32]);
wire tmp_7_33;
assign tmp_7_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_7_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_7_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_7_V_read[33]);
wire tmp_7_34;
assign tmp_7_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_7_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_7_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_7_V_read[34]);
wire tmp_7_35;
assign tmp_7_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_7_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_7_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_7_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_7_V_read[35]);
wire tmp_7_36;
assign tmp_7_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_7_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_7_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_7_V_read[36]);
wire tmp_7_37;
assign tmp_7_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_7_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_7_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_7_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_7_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_7_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_7_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_7_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_7_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_7_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_7_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_7_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_7_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_7_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_7_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_7_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_7_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_7_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_7_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_7_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_7_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_7_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_7_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_7_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_7_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_7_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_7_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_7_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_7_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_7_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_7_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_7_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_7_V_read[37]);
wire tmp_7_38;
assign tmp_7_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_7_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_7_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_7_V_read[38]);
wire tmp_7_40;
assign tmp_7_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_7_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_7_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_7_V_read[40]);
wire tmp_7_41;
assign tmp_7_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_7_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_7_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_7_V_read[41]);
wire tmp_7_42;
assign tmp_7_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_7_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_7_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_7_V_read[42]);
wire tmp_7_43;
assign tmp_7_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_7_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_7_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_7_V_read[43]);
wire tmp_7_44;
assign tmp_7_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_7_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_7_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_7_V_read[44]);
wire tmp_7_45;
assign tmp_7_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_7_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_7_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_7_V_read[45]);
wire tmp_7_46;
assign tmp_7_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_7_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_7_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_7_V_read[46]);
wire tmp_7_47;
assign tmp_7_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_7_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_7_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_7_V_read[47]);
wire tmp_7_48;
assign tmp_7_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_7_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_7_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_7_V_read[48]);
wire tmp_7_49;
assign tmp_7_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_7_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_7_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_7_V_read[49]);
wire tmp_7_50;
assign tmp_7_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_7_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_7_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_7_V_read[50]);
wire tmp_7_51;
assign tmp_7_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_7_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_7_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_7_V_read[51]);
wire tmp_7_52;
assign tmp_7_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_7_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_7_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_7_V_read[52]);
wire tmp_7_53;
assign tmp_7_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_7_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_7_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_7_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_7_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_7_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_7_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_7_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_7_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_7_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_7_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_7_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_7_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_7_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_7_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_7_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_7_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_7_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_7_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_7_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_7_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_7_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_7_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_7_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_7_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_7_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_7_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_7_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_7_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_7_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_7_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_7_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_7_V_read[53]);
wire tmp_7_54;
assign tmp_7_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_7_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_7_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_7_V_read[54]);
wire tmp_7_55;
assign tmp_7_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_7_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_7_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_7_V_read[55]);
wire tmp_7_56;
assign tmp_7_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_7_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_7_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_7_V_read[56]);
wire tmp_7_57;
assign tmp_7_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_7_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_7_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_7_V_read[57]);
wire tmp_7_58;
assign tmp_7_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_7_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_7_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_7_V_read[58]);
wire tmp_7_60;
assign tmp_7_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_7_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_7_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_7_V_read[60]);
wire tmp_7_61;
assign tmp_7_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_7_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_7_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_7_V_read[61]);
wire tmp_7_62;
assign tmp_7_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_7_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_7_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_7_V_read[62]);
wire tmp_7_64;
assign tmp_7_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_7_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_7_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_7_V_read[64]);
wire tmp_7_65;
assign tmp_7_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_7_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_7_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_7_V_read[65]);
wire tmp_7_66;
assign tmp_7_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_7_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_7_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_7_V_read[66]);
wire tmp_7_67;
assign tmp_7_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_7_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_7_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_7_V_read[67]);
wire tmp_7_68;
assign tmp_7_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_7_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_7_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_7_V_read[68]);
wire tmp_7_69;
assign tmp_7_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_7_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_7_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_7_V_read[69]);
wire tmp_7_70;
assign tmp_7_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_7_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_7_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_7_V_read[70]);
assign ap_return_7 = {tmp_7_0,tmp_7_1,tmp_7_2,tmp_7_3,tmp_7_4,tmp_7_5,tmp_7_6,tmp_7_7,1'b0,tmp_7_9,tmp_7_10,1'b0,tmp_7_12,tmp_7_13,tmp_7_14,tmp_7_15,tmp_7_16,tmp_7_17,tmp_7_18,tmp_7_19,tmp_7_20,tmp_7_21,tmp_7_22,tmp_7_23,tmp_7_24,1'b0,tmp_7_26,tmp_7_27,tmp_7_28,tmp_7_29,tmp_7_30,tmp_7_31,tmp_7_32,tmp_7_33,tmp_7_34,tmp_7_35,tmp_7_36,tmp_7_37,tmp_7_38,1'b0,tmp_7_40,tmp_7_41,tmp_7_42,tmp_7_43,tmp_7_44,tmp_7_45,tmp_7_46,tmp_7_47,tmp_7_48,tmp_7_49,tmp_7_50,tmp_7_51,tmp_7_52,tmp_7_53,tmp_7_54,tmp_7_55,tmp_7_56,tmp_7_57,tmp_7_58,1'b0,tmp_7_60,tmp_7_61,tmp_7_62,1'b0,tmp_7_64,tmp_7_65,tmp_7_66,tmp_7_67,tmp_7_68,tmp_7_69,tmp_7_70,1'b0};
wire tmp_8_0;
assign tmp_8_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_8_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_8_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_8_V_read[0]);
wire tmp_8_1;
assign tmp_8_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_8_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_8_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_8_V_read[1]);
wire tmp_8_2;
assign tmp_8_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_8_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_8_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_8_V_read[2]);
wire tmp_8_3;
assign tmp_8_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_8_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_8_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_8_V_read[3]);
wire tmp_8_5;
assign tmp_8_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_8_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_8_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_8_V_read[5]);
wire tmp_8_6;
assign tmp_8_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_8_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_8_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_8_V_read[6]);
wire tmp_8_8;
assign tmp_8_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_8_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_8_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_8_V_read[8]);
wire tmp_8_9;
assign tmp_8_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_8_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_8_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_8_V_read[9]);
wire tmp_8_10;
assign tmp_8_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_8_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_8_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_8_V_read[10]);
wire tmp_8_11;
assign tmp_8_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_8_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_8_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_8_V_read[11]);
wire tmp_8_12;
assign tmp_8_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_8_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_8_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_8_V_read[12]);
wire tmp_8_13;
assign tmp_8_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_8_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_8_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_8_V_read[13]);
wire tmp_8_14;
assign tmp_8_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_8_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_8_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_8_V_read[14]);
wire tmp_8_16;
assign tmp_8_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_8_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_8_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_8_V_read[16]);
wire tmp_8_17;
assign tmp_8_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_8_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_8_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_8_V_read[17]);
wire tmp_8_18;
assign tmp_8_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_8_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_8_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_8_V_read[18]);
wire tmp_8_19;
assign tmp_8_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_8_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_8_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_8_V_read[19]);
wire tmp_8_20;
assign tmp_8_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_8_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_8_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_8_V_read[20]);
wire tmp_8_21;
assign tmp_8_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_8_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_8_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_8_V_read[21]);
wire tmp_8_22;
assign tmp_8_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_8_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_8_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_8_V_read[22]);
wire tmp_8_23;
assign tmp_8_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_8_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_8_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_8_V_read[23]);
wire tmp_8_24;
assign tmp_8_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_8_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_8_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_8_V_read[24]);
wire tmp_8_25;
assign tmp_8_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_8_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_8_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_8_V_read[25]);
wire tmp_8_26;
assign tmp_8_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_8_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_8_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_8_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_8_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_8_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_8_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_8_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_8_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_8_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_8_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_8_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_8_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_8_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_8_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_8_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_8_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_8_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_8_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_8_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_8_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_8_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_8_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_8_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_8_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_8_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_8_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_8_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_8_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_8_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_8_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_8_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_8_V_read[26]);
wire tmp_8_27;
assign tmp_8_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_8_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_8_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_8_V_read[27]);
wire tmp_8_28;
assign tmp_8_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_8_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_8_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_8_V_read[28]);
wire tmp_8_29;
assign tmp_8_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_8_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_8_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_8_V_read[29]);
wire tmp_8_30;
assign tmp_8_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_8_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_8_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_8_V_read[30]);
wire tmp_8_32;
assign tmp_8_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_8_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_8_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_8_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_8_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_8_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_8_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_8_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_8_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_8_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_8_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_8_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_8_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_8_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_8_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_8_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_8_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_8_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_8_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_8_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_8_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_8_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_8_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_8_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_8_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_8_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_8_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_8_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_8_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_8_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_8_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_8_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_8_V_read[32]);
wire tmp_8_33;
assign tmp_8_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_8_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_8_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_8_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_8_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_8_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_8_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_8_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_8_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_8_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_8_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_8_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_8_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_8_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_8_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_8_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_8_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_8_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_8_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_8_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_8_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_8_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_8_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_8_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_8_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_8_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_8_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_8_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_8_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_8_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_8_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_8_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_8_V_read[33]);
wire tmp_8_34;
assign tmp_8_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_8_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_8_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_8_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_8_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_8_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_8_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_8_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_8_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_8_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_8_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_8_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_8_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_8_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_8_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_8_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_8_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_8_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_8_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_8_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_8_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_8_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_8_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_8_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_8_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_8_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_8_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_8_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_8_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_8_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_8_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_8_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_8_V_read[34]);
wire tmp_8_35;
assign tmp_8_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_8_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_8_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_8_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_8_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_8_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_8_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_8_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_8_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_8_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_8_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_8_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_8_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_8_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_8_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_8_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_8_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_8_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_8_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_8_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_8_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_8_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_8_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_8_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_8_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_8_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_8_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_8_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_8_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_8_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_8_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_8_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_8_V_read[35]);
wire tmp_8_36;
assign tmp_8_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_8_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_8_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_8_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_8_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_8_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_8_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_8_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_8_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_8_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_8_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_8_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_8_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_8_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_8_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_8_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_8_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_8_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_8_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_8_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_8_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_8_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_8_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_8_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_8_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_8_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_8_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_8_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_8_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_8_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_8_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_8_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_8_V_read[36]);
wire tmp_8_37;
assign tmp_8_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_8_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_8_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_8_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_8_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_8_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_8_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_8_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_8_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_8_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_8_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_8_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_8_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_8_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_8_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_8_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_8_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_8_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_8_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_8_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_8_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_8_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_8_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_8_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_8_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_8_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_8_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_8_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_8_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_8_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_8_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_8_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_8_V_read[37]);
wire tmp_8_38;
assign tmp_8_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_8_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_8_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_8_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_8_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_8_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_8_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_8_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_8_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_8_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_8_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_8_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_8_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_8_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_8_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_8_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_8_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_8_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_8_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_8_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_8_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_8_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_8_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_8_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_8_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_8_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_8_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_8_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_8_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_8_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_8_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_8_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_8_V_read[38]);
wire tmp_8_39;
assign tmp_8_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_8_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_8_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_8_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_8_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_8_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_8_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_8_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_8_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_8_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_8_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_8_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_8_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_8_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_8_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_8_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_8_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_8_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_8_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_8_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_8_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_8_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_8_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_8_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_8_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_8_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_8_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_8_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_8_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_8_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_8_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_8_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_8_V_read[39]);
wire tmp_8_40;
assign tmp_8_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_8_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_8_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_8_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_8_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_8_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_8_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_8_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_8_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_8_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_8_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_8_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_8_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_8_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_8_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_8_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_8_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_8_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_8_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_8_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_8_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_8_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_8_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_8_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_8_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_8_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_8_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_8_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_8_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_8_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_8_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_8_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_8_V_read[40]);
wire tmp_8_42;
assign tmp_8_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_8_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_8_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_8_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_8_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_8_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_8_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_8_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_8_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_8_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_8_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_8_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_8_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_8_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_8_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_8_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_8_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_8_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_8_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_8_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_8_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_8_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_8_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_8_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_8_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_8_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_8_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_8_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_8_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_8_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_8_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_8_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_8_V_read[42]);
wire tmp_8_43;
assign tmp_8_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_8_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_8_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_8_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_8_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_8_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_8_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_8_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_8_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_8_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_8_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_8_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_8_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_8_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_8_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_8_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_8_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_8_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_8_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_8_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_8_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_8_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_8_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_8_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_8_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_8_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_8_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_8_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_8_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_8_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_8_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_8_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_8_V_read[43]);
wire tmp_8_44;
assign tmp_8_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_8_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_8_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_8_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_8_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_8_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_8_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_8_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_8_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_8_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_8_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_8_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_8_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_8_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_8_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_8_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_8_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_8_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_8_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_8_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_8_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_8_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_8_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_8_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_8_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_8_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_8_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_8_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_8_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_8_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_8_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_8_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_8_V_read[44]);
wire tmp_8_45;
assign tmp_8_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_8_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_8_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_8_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_8_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_8_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_8_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_8_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_8_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_8_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_8_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_8_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_8_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_8_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_8_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_8_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_8_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_8_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_8_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_8_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_8_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_8_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_8_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_8_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_8_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_8_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_8_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_8_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_8_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_8_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_8_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_8_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_8_V_read[45]);
wire tmp_8_46;
assign tmp_8_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_8_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_8_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_8_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_8_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_8_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_8_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_8_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_8_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_8_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_8_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_8_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_8_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_8_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_8_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_8_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_8_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_8_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_8_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_8_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_8_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_8_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_8_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_8_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_8_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_8_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_8_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_8_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_8_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_8_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_8_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_8_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_8_V_read[46]);
wire tmp_8_47;
assign tmp_8_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_8_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_8_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_8_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_8_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_8_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_8_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_8_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_8_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_8_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_8_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_8_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_8_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_8_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_8_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_8_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_8_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_8_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_8_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_8_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_8_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_8_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_8_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_8_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_8_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_8_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_8_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_8_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_8_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_8_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_8_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_8_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_8_V_read[47]);
wire tmp_8_48;
assign tmp_8_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_8_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_8_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_8_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_8_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_8_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_8_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_8_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_8_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_8_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_8_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_8_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_8_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_8_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_8_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_8_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_8_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_8_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_8_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_8_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_8_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_8_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_8_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_8_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_8_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_8_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_8_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_8_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_8_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_8_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_8_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_8_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_8_V_read[48]);
wire tmp_8_49;
assign tmp_8_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_8_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_8_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_8_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_8_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_8_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_8_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_8_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_8_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_8_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_8_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_8_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_8_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_8_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_8_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_8_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_8_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_8_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_8_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_8_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_8_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_8_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_8_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_8_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_8_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_8_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_8_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_8_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_8_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_8_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_8_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_8_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_8_V_read[49]);
wire tmp_8_50;
assign tmp_8_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_8_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_8_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_8_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_8_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_8_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_8_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_8_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_8_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_8_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_8_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_8_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_8_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_8_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_8_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_8_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_8_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_8_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_8_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_8_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_8_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_8_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_8_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_8_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_8_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_8_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_8_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_8_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_8_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_8_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_8_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_8_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_8_V_read[50]);
wire tmp_8_51;
assign tmp_8_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_8_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_8_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_8_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_8_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_8_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_8_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_8_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_8_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_8_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_8_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_8_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_8_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_8_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_8_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_8_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_8_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_8_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_8_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_8_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_8_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_8_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_8_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_8_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_8_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_8_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_8_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_8_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_8_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_8_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_8_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_8_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_8_V_read[51]);
wire tmp_8_52;
assign tmp_8_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_8_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_8_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_8_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_8_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_8_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_8_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_8_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_8_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_8_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_8_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_8_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_8_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_8_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_8_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_8_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_8_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_8_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_8_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_8_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_8_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_8_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_8_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_8_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_8_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_8_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_8_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_8_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_8_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_8_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_8_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_8_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_8_V_read[52]);
wire tmp_8_53;
assign tmp_8_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_8_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_8_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_8_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_8_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_8_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_8_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_8_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_8_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_8_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_8_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_8_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_8_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_8_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_8_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_8_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_8_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_8_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_8_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_8_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_8_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_8_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_8_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_8_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_8_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_8_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_8_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_8_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_8_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_8_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_8_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_8_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_8_V_read[53]);
wire tmp_8_54;
assign tmp_8_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_8_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_8_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_8_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_8_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_8_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_8_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_8_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_8_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_8_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_8_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_8_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_8_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_8_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_8_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_8_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_8_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_8_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_8_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_8_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_8_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_8_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_8_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_8_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_8_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_8_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_8_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_8_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_8_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_8_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_8_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_8_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_8_V_read[54]);
wire tmp_8_55;
assign tmp_8_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_8_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_8_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_8_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_8_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_8_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_8_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_8_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_8_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_8_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_8_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_8_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_8_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_8_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_8_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_8_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_8_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_8_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_8_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_8_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_8_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_8_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_8_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_8_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_8_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_8_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_8_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_8_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_8_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_8_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_8_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_8_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_8_V_read[55]);
wire tmp_8_56;
assign tmp_8_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_8_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_8_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_8_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_8_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_8_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_8_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_8_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_8_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_8_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_8_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_8_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_8_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_8_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_8_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_8_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_8_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_8_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_8_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_8_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_8_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_8_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_8_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_8_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_8_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_8_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_8_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_8_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_8_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_8_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_8_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_8_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_8_V_read[56]);
wire tmp_8_57;
assign tmp_8_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_8_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_8_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_8_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_8_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_8_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_8_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_8_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_8_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_8_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_8_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_8_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_8_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_8_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_8_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_8_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_8_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_8_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_8_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_8_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_8_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_8_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_8_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_8_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_8_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_8_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_8_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_8_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_8_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_8_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_8_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_8_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_8_V_read[57]);
wire tmp_8_58;
assign tmp_8_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_8_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_8_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_8_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_8_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_8_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_8_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_8_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_8_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_8_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_8_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_8_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_8_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_8_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_8_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_8_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_8_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_8_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_8_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_8_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_8_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_8_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_8_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_8_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_8_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_8_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_8_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_8_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_8_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_8_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_8_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_8_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_8_V_read[58]);
wire tmp_8_59;
assign tmp_8_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_8_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_8_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_8_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_8_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_8_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_8_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_8_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_8_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_8_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_8_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_8_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_8_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_8_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_8_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_8_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_8_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_8_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_8_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_8_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_8_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_8_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_8_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_8_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_8_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_8_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_8_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_8_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_8_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_8_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_8_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_8_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_8_V_read[59]);
wire tmp_8_60;
assign tmp_8_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_8_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_8_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_8_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_8_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_8_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_8_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_8_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_8_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_8_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_8_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_8_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_8_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_8_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_8_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_8_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_8_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_8_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_8_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_8_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_8_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_8_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_8_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_8_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_8_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_8_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_8_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_8_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_8_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_8_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_8_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_8_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_8_V_read[60]);
wire tmp_8_61;
assign tmp_8_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_8_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_8_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_8_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_8_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_8_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_8_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_8_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_8_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_8_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_8_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_8_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_8_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_8_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_8_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_8_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_8_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_8_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_8_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_8_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_8_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_8_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_8_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_8_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_8_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_8_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_8_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_8_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_8_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_8_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_8_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_8_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_8_V_read[61]);
wire tmp_8_62;
assign tmp_8_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_8_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_8_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_8_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_8_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_8_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_8_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_8_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_8_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_8_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_8_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_8_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_8_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_8_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_8_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_8_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_8_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_8_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_8_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_8_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_8_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_8_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_8_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_8_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_8_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_8_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_8_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_8_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_8_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_8_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_8_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_8_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_8_V_read[62]);
wire tmp_8_65;
assign tmp_8_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_8_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_8_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_8_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_8_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_8_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_8_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_8_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_8_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_8_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_8_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_8_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_8_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_8_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_8_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_8_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_8_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_8_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_8_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_8_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_8_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_8_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_8_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_8_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_8_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_8_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_8_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_8_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_8_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_8_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_8_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_8_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_8_V_read[65]);
wire tmp_8_66;
assign tmp_8_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_8_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_8_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_8_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_8_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_8_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_8_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_8_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_8_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_8_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_8_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_8_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_8_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_8_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_8_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_8_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_8_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_8_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_8_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_8_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_8_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_8_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_8_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_8_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_8_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_8_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_8_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_8_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_8_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_8_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_8_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_8_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_8_V_read[66]);
wire tmp_8_67;
assign tmp_8_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_8_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_8_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_8_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_8_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_8_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_8_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_8_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_8_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_8_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_8_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_8_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_8_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_8_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_8_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_8_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_8_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_8_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_8_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_8_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_8_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_8_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_8_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_8_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_8_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_8_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_8_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_8_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_8_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_8_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_8_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_8_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_8_V_read[67]);
wire tmp_8_69;
assign tmp_8_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_8_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_8_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_8_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_8_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_8_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_8_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_8_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_8_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_8_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_8_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_8_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_8_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_8_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_8_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_8_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_8_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_8_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_8_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_8_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_8_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_8_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_8_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_8_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_8_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_8_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_8_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_8_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_8_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_8_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_8_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_8_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_8_V_read[69]);
wire tmp_8_70;
assign tmp_8_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_8_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_8_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_8_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_8_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_8_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_8_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_8_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_8_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_8_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_8_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_8_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_8_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_8_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_8_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_8_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_8_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_8_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_8_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_8_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_8_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_8_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_8_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_8_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_8_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_8_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_8_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_8_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_8_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_8_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_8_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_8_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_8_V_read[70]);
wire tmp_8_71;
assign tmp_8_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_8_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_8_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_8_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_8_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_8_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_8_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_8_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_8_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_8_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_8_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_8_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_8_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_8_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_8_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_8_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_8_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_8_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_8_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_8_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_8_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_8_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_8_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_8_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_8_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_8_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_8_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_8_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_8_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_8_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_8_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_8_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_8_V_read[71]);
assign ap_return_8 = {tmp_8_0,tmp_8_1,tmp_8_2,tmp_8_3,1'b0,tmp_8_5,tmp_8_6,1'b0,tmp_8_8,tmp_8_9,tmp_8_10,tmp_8_11,tmp_8_12,tmp_8_13,tmp_8_14,1'b0,tmp_8_16,tmp_8_17,tmp_8_18,tmp_8_19,tmp_8_20,tmp_8_21,tmp_8_22,tmp_8_23,tmp_8_24,tmp_8_25,tmp_8_26,tmp_8_27,tmp_8_28,tmp_8_29,tmp_8_30,1'b0,tmp_8_32,tmp_8_33,tmp_8_34,tmp_8_35,tmp_8_36,tmp_8_37,tmp_8_38,tmp_8_39,tmp_8_40,1'b0,tmp_8_42,tmp_8_43,tmp_8_44,tmp_8_45,tmp_8_46,tmp_8_47,tmp_8_48,tmp_8_49,tmp_8_50,tmp_8_51,tmp_8_52,tmp_8_53,tmp_8_54,tmp_8_55,tmp_8_56,tmp_8_57,tmp_8_58,tmp_8_59,tmp_8_60,tmp_8_61,tmp_8_62,1'b0,1'b0,tmp_8_65,tmp_8_66,tmp_8_67,1'b0,tmp_8_69,tmp_8_70,tmp_8_71};
wire tmp_9_0;
assign tmp_9_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_9_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_9_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_9_V_read[0]);
wire tmp_9_1;
assign tmp_9_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_9_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_9_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_9_V_read[1]);
wire tmp_9_2;
assign tmp_9_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_9_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_9_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_9_V_read[2]);
wire tmp_9_3;
assign tmp_9_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_9_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_9_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_9_V_read[3]);
wire tmp_9_4;
assign tmp_9_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_9_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_9_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_9_V_read[4]);
wire tmp_9_5;
assign tmp_9_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_9_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_9_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_9_V_read[5]);
wire tmp_9_7;
assign tmp_9_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_9_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_9_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_9_V_read[7]);
wire tmp_9_8;
assign tmp_9_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_9_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_9_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_9_V_read[8]);
wire tmp_9_9;
assign tmp_9_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_9_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_9_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_9_V_read[9]);
wire tmp_9_10;
assign tmp_9_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_9_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_9_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_9_V_read[10]);
wire tmp_9_11;
assign tmp_9_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_9_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_9_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_9_V_read[11]);
wire tmp_9_12;
assign tmp_9_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_9_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_9_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_9_V_read[12]);
wire tmp_9_13;
assign tmp_9_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_9_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_9_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_9_V_read[13]);
wire tmp_9_14;
assign tmp_9_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_9_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_9_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_9_V_read[14]);
wire tmp_9_15;
assign tmp_9_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_9_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_9_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_9_V_read[15]);
wire tmp_9_16;
assign tmp_9_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_9_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_9_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_9_V_read[16]);
wire tmp_9_17;
assign tmp_9_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_9_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_9_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_9_V_read[17]);
wire tmp_9_18;
assign tmp_9_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_9_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_9_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_9_V_read[18]);
wire tmp_9_19;
assign tmp_9_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_9_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_9_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_9_V_read[19]);
wire tmp_9_20;
assign tmp_9_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_9_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_9_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_9_V_read[20]);
wire tmp_9_21;
assign tmp_9_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_9_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_9_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_9_V_read[21]);
wire tmp_9_22;
assign tmp_9_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_9_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_9_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_9_V_read[22]);
wire tmp_9_23;
assign tmp_9_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_9_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_9_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_9_V_read[23]);
wire tmp_9_24;
assign tmp_9_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_9_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_9_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_9_V_read[24]);
wire tmp_9_25;
assign tmp_9_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_9_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_9_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_9_V_read[25]);
wire tmp_9_26;
assign tmp_9_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_9_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_9_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_9_V_read[26]);
wire tmp_9_27;
assign tmp_9_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_9_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_9_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_9_V_read[27]);
wire tmp_9_28;
assign tmp_9_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_9_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_9_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_9_V_read[28]);
wire tmp_9_29;
assign tmp_9_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_9_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_9_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_9_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_9_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_9_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_9_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_9_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_9_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_9_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_9_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_9_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_9_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_9_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_9_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_9_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_9_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_9_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_9_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_9_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_9_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_9_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_9_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_9_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_9_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_9_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_9_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_9_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_9_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_9_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_9_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_9_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_9_V_read[29]);
wire tmp_9_31;
assign tmp_9_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_9_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_9_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_9_V_read[31]);
wire tmp_9_33;
assign tmp_9_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_9_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_9_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_9_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_9_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_9_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_9_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_9_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_9_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_9_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_9_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_9_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_9_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_9_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_9_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_9_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_9_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_9_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_9_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_9_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_9_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_9_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_9_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_9_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_9_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_9_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_9_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_9_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_9_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_9_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_9_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_9_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_9_V_read[33]);
wire tmp_9_34;
assign tmp_9_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_9_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_9_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_9_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_9_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_9_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_9_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_9_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_9_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_9_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_9_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_9_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_9_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_9_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_9_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_9_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_9_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_9_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_9_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_9_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_9_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_9_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_9_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_9_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_9_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_9_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_9_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_9_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_9_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_9_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_9_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_9_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_9_V_read[34]);
wire tmp_9_35;
assign tmp_9_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_9_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_9_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_9_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_9_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_9_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_9_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_9_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_9_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_9_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_9_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_9_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_9_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_9_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_9_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_9_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_9_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_9_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_9_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_9_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_9_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_9_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_9_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_9_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_9_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_9_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_9_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_9_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_9_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_9_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_9_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_9_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_9_V_read[35]);
wire tmp_9_37;
assign tmp_9_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_9_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_9_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_9_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_9_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_9_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_9_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_9_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_9_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_9_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_9_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_9_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_9_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_9_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_9_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_9_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_9_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_9_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_9_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_9_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_9_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_9_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_9_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_9_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_9_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_9_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_9_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_9_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_9_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_9_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_9_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_9_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_9_V_read[37]);
wire tmp_9_38;
assign tmp_9_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_9_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_9_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_9_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_9_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_9_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_9_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_9_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_9_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_9_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_9_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_9_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_9_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_9_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_9_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_9_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_9_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_9_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_9_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_9_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_9_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_9_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_9_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_9_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_9_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_9_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_9_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_9_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_9_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_9_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_9_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_9_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_9_V_read[38]);
wire tmp_9_40;
assign tmp_9_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_9_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_9_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_9_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_9_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_9_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_9_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_9_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_9_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_9_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_9_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_9_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_9_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_9_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_9_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_9_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_9_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_9_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_9_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_9_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_9_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_9_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_9_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_9_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_9_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_9_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_9_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_9_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_9_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_9_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_9_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_9_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_9_V_read[40]);
wire tmp_9_41;
assign tmp_9_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_9_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_9_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_9_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_9_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_9_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_9_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_9_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_9_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_9_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_9_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_9_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_9_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_9_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_9_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_9_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_9_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_9_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_9_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_9_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_9_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_9_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_9_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_9_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_9_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_9_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_9_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_9_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_9_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_9_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_9_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_9_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_9_V_read[41]);
wire tmp_9_42;
assign tmp_9_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_9_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_9_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_9_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_9_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_9_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_9_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_9_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_9_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_9_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_9_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_9_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_9_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_9_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_9_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_9_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_9_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_9_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_9_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_9_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_9_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_9_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_9_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_9_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_9_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_9_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_9_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_9_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_9_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_9_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_9_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_9_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_9_V_read[42]);
wire tmp_9_43;
assign tmp_9_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_9_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_9_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_9_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_9_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_9_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_9_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_9_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_9_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_9_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_9_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_9_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_9_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_9_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_9_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_9_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_9_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_9_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_9_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_9_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_9_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_9_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_9_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_9_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_9_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_9_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_9_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_9_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_9_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_9_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_9_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_9_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_9_V_read[43]);
wire tmp_9_44;
assign tmp_9_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_9_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_9_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_9_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_9_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_9_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_9_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_9_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_9_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_9_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_9_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_9_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_9_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_9_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_9_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_9_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_9_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_9_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_9_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_9_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_9_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_9_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_9_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_9_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_9_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_9_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_9_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_9_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_9_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_9_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_9_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_9_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_9_V_read[44]);
wire tmp_9_45;
assign tmp_9_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_9_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_9_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_9_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_9_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_9_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_9_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_9_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_9_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_9_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_9_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_9_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_9_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_9_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_9_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_9_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_9_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_9_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_9_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_9_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_9_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_9_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_9_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_9_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_9_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_9_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_9_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_9_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_9_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_9_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_9_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_9_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_9_V_read[45]);
wire tmp_9_46;
assign tmp_9_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_9_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_9_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_9_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_9_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_9_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_9_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_9_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_9_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_9_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_9_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_9_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_9_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_9_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_9_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_9_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_9_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_9_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_9_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_9_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_9_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_9_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_9_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_9_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_9_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_9_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_9_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_9_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_9_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_9_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_9_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_9_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_9_V_read[46]);
wire tmp_9_47;
assign tmp_9_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_9_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_9_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_9_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_9_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_9_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_9_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_9_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_9_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_9_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_9_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_9_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_9_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_9_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_9_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_9_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_9_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_9_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_9_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_9_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_9_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_9_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_9_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_9_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_9_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_9_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_9_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_9_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_9_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_9_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_9_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_9_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_9_V_read[47]);
wire tmp_9_48;
assign tmp_9_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_9_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_9_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_9_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_9_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_9_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_9_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_9_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_9_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_9_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_9_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_9_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_9_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_9_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_9_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_9_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_9_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_9_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_9_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_9_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_9_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_9_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_9_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_9_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_9_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_9_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_9_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_9_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_9_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_9_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_9_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_9_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_9_V_read[48]);
wire tmp_9_49;
assign tmp_9_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_9_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_9_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_9_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_9_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_9_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_9_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_9_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_9_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_9_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_9_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_9_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_9_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_9_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_9_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_9_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_9_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_9_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_9_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_9_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_9_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_9_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_9_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_9_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_9_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_9_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_9_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_9_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_9_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_9_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_9_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_9_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_9_V_read[49]);
wire tmp_9_50;
assign tmp_9_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_9_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_9_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_9_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_9_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_9_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_9_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_9_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_9_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_9_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_9_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_9_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_9_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_9_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_9_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_9_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_9_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_9_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_9_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_9_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_9_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_9_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_9_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_9_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_9_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_9_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_9_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_9_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_9_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_9_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_9_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_9_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_9_V_read[50]);
wire tmp_9_51;
assign tmp_9_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_9_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_9_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_9_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_9_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_9_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_9_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_9_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_9_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_9_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_9_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_9_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_9_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_9_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_9_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_9_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_9_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_9_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_9_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_9_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_9_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_9_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_9_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_9_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_9_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_9_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_9_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_9_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_9_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_9_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_9_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_9_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_9_V_read[51]);
wire tmp_9_52;
assign tmp_9_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_9_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_9_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_9_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_9_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_9_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_9_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_9_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_9_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_9_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_9_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_9_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_9_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_9_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_9_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_9_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_9_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_9_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_9_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_9_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_9_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_9_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_9_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_9_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_9_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_9_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_9_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_9_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_9_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_9_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_9_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_9_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_9_V_read[52]);
wire tmp_9_53;
assign tmp_9_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_9_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_9_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_9_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_9_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_9_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_9_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_9_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_9_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_9_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_9_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_9_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_9_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_9_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_9_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_9_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_9_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_9_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_9_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_9_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_9_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_9_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_9_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_9_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_9_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_9_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_9_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_9_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_9_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_9_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_9_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_9_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_9_V_read[53]);
wire tmp_9_54;
assign tmp_9_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_9_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_9_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_9_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_9_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_9_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_9_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_9_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_9_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_9_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_9_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_9_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_9_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_9_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_9_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_9_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_9_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_9_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_9_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_9_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_9_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_9_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_9_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_9_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_9_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_9_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_9_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_9_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_9_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_9_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_9_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_9_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_9_V_read[54]);
wire tmp_9_55;
assign tmp_9_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_9_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_9_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_9_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_9_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_9_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_9_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_9_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_9_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_9_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_9_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_9_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_9_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_9_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_9_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_9_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_9_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_9_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_9_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_9_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_9_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_9_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_9_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_9_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_9_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_9_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_9_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_9_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_9_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_9_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_9_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_9_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_9_V_read[55]);
wire tmp_9_56;
assign tmp_9_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_9_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_9_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_9_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_9_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_9_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_9_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_9_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_9_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_9_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_9_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_9_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_9_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_9_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_9_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_9_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_9_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_9_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_9_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_9_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_9_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_9_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_9_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_9_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_9_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_9_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_9_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_9_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_9_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_9_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_9_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_9_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_9_V_read[56]);
wire tmp_9_57;
assign tmp_9_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_9_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_9_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_9_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_9_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_9_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_9_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_9_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_9_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_9_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_9_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_9_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_9_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_9_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_9_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_9_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_9_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_9_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_9_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_9_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_9_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_9_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_9_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_9_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_9_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_9_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_9_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_9_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_9_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_9_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_9_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_9_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_9_V_read[57]);
wire tmp_9_58;
assign tmp_9_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_9_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_9_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_9_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_9_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_9_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_9_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_9_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_9_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_9_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_9_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_9_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_9_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_9_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_9_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_9_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_9_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_9_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_9_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_9_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_9_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_9_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_9_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_9_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_9_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_9_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_9_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_9_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_9_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_9_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_9_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_9_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_9_V_read[58]);
wire tmp_9_59;
assign tmp_9_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_9_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_9_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_9_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_9_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_9_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_9_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_9_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_9_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_9_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_9_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_9_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_9_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_9_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_9_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_9_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_9_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_9_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_9_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_9_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_9_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_9_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_9_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_9_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_9_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_9_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_9_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_9_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_9_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_9_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_9_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_9_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_9_V_read[59]);
wire tmp_9_60;
assign tmp_9_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_9_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_9_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_9_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_9_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_9_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_9_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_9_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_9_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_9_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_9_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_9_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_9_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_9_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_9_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_9_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_9_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_9_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_9_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_9_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_9_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_9_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_9_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_9_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_9_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_9_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_9_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_9_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_9_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_9_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_9_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_9_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_9_V_read[60]);
wire tmp_9_61;
assign tmp_9_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_9_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_9_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_9_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_9_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_9_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_9_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_9_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_9_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_9_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_9_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_9_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_9_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_9_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_9_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_9_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_9_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_9_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_9_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_9_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_9_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_9_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_9_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_9_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_9_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_9_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_9_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_9_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_9_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_9_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_9_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_9_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_9_V_read[61]);
wire tmp_9_62;
assign tmp_9_62 = (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_9_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_9_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_9_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_9_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_9_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_9_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_9_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_9_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_9_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_9_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_9_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_9_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_9_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_9_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_9_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_9_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_9_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_9_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_9_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_9_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_9_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_9_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_9_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_9_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_9_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_9_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_9_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_9_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_9_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_9_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_9_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_9_V_read[62]);
wire tmp_9_63;
assign tmp_9_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_9_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_9_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_9_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_9_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_9_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_9_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_9_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_9_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_9_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_9_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_9_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_9_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_9_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_9_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_9_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_9_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_9_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_9_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_9_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_9_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_9_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_9_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_9_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_9_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_9_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_9_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_9_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_9_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_9_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_9_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_9_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_9_V_read[63]);
wire tmp_9_64;
assign tmp_9_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_9_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_9_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_9_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_9_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_9_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_9_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_9_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_9_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_9_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_9_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_9_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_9_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_9_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_9_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_9_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_9_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_9_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_9_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_9_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_9_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_9_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_9_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_9_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_9_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_9_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_9_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_9_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_9_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_9_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_9_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_9_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_9_V_read[64]);
wire tmp_9_65;
assign tmp_9_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_9_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_9_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_9_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_9_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_9_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_9_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_9_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_9_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_9_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_9_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_9_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_9_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_9_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_9_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_9_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_9_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_9_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_9_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_9_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_9_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_9_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_9_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_9_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_9_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_9_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_9_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_9_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_9_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_9_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_9_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_9_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_9_V_read[65]);
wire tmp_9_67;
assign tmp_9_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_9_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_9_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_9_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_9_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_9_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_9_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_9_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_9_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_9_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_9_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_9_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_9_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_9_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_9_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_9_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_9_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_9_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_9_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_9_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_9_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_9_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_9_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_9_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_9_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_9_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_9_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_9_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_9_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_9_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_9_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_9_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_9_V_read[67]);
wire tmp_9_68;
assign tmp_9_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_9_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_9_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_9_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_9_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_9_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_9_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_9_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_9_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_9_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_9_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_9_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_9_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_9_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_9_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_9_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_9_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_9_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_9_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_9_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_9_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_9_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_9_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_9_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_9_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_9_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_9_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_9_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_9_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_9_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_9_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_9_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_9_V_read[68]);
wire tmp_9_69;
assign tmp_9_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_9_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_9_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_9_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_9_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_9_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_9_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_9_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_9_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_9_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_9_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_9_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_9_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_9_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_9_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_9_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_9_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_9_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_9_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_9_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_9_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_9_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_9_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_9_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_9_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_9_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_9_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_9_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_9_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_9_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_9_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_9_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_9_V_read[69]);
wire tmp_9_70;
assign tmp_9_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_9_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_9_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_9_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_9_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_9_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_9_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_9_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_9_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_9_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_9_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_9_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_9_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_9_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_9_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_9_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_9_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_9_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_9_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_9_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_9_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_9_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_9_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_9_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_9_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_9_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_9_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_9_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_9_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_9_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_9_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_9_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_9_V_read[70]);
wire tmp_9_71;
assign tmp_9_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_9_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_9_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_9_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_9_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_9_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_9_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_9_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_9_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_9_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_9_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_9_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_9_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_9_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_9_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_9_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_9_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_9_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_9_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_9_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_9_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_9_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_9_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_9_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_9_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_9_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_9_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_9_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_9_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_9_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_9_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_9_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_9_V_read[71]);
assign ap_return_9 = {tmp_9_0,tmp_9_1,tmp_9_2,tmp_9_3,tmp_9_4,tmp_9_5,1'b0,tmp_9_7,tmp_9_8,tmp_9_9,tmp_9_10,tmp_9_11,tmp_9_12,tmp_9_13,tmp_9_14,tmp_9_15,tmp_9_16,tmp_9_17,tmp_9_18,tmp_9_19,tmp_9_20,tmp_9_21,tmp_9_22,tmp_9_23,tmp_9_24,tmp_9_25,tmp_9_26,tmp_9_27,tmp_9_28,tmp_9_29,1'b0,tmp_9_31,1'b0,tmp_9_33,tmp_9_34,tmp_9_35,1'b0,tmp_9_37,tmp_9_38,1'b0,tmp_9_40,tmp_9_41,tmp_9_42,tmp_9_43,tmp_9_44,tmp_9_45,tmp_9_46,tmp_9_47,tmp_9_48,tmp_9_49,tmp_9_50,tmp_9_51,tmp_9_52,tmp_9_53,tmp_9_54,tmp_9_55,tmp_9_56,tmp_9_57,tmp_9_58,tmp_9_59,tmp_9_60,tmp_9_61,tmp_9_62,tmp_9_63,tmp_9_64,tmp_9_65,1'b0,tmp_9_67,tmp_9_68,tmp_9_69,tmp_9_70,tmp_9_71};
wire tmp_10_0;
assign tmp_10_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_10_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_10_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_10_V_read[0]);
wire tmp_10_1;
assign tmp_10_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_10_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_10_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_10_V_read[1]);
wire tmp_10_2;
assign tmp_10_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_10_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_10_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_10_V_read[2]);
wire tmp_10_3;
assign tmp_10_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_10_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_10_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_10_V_read[3]);
wire tmp_10_4;
assign tmp_10_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_10_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_10_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_10_V_read[4]);
wire tmp_10_5;
assign tmp_10_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_10_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_10_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_10_V_read[5]);
wire tmp_10_6;
assign tmp_10_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_10_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_10_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_10_V_read[6]);
wire tmp_10_7;
assign tmp_10_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_10_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_10_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_10_V_read[7]);
wire tmp_10_8;
assign tmp_10_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_10_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_10_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_10_V_read[8]);
wire tmp_10_9;
assign tmp_10_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_10_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_10_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_10_V_read[9]);
wire tmp_10_10;
assign tmp_10_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_10_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_10_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_10_V_read[10]);
wire tmp_10_11;
assign tmp_10_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_10_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_10_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_10_V_read[11]);
wire tmp_10_12;
assign tmp_10_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_10_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_10_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_10_V_read[12]);
wire tmp_10_13;
assign tmp_10_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_10_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_10_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_10_V_read[13]);
wire tmp_10_14;
assign tmp_10_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_10_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_10_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_10_V_read[14]);
wire tmp_10_15;
assign tmp_10_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_10_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_10_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_10_V_read[15]);
wire tmp_10_16;
assign tmp_10_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_10_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_10_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_10_V_read[16]);
wire tmp_10_17;
assign tmp_10_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_10_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_10_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_10_V_read[17]);
wire tmp_10_19;
assign tmp_10_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_10_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_10_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_10_V_read[19]);
wire tmp_10_20;
assign tmp_10_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_10_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_10_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_10_V_read[20]);
wire tmp_10_21;
assign tmp_10_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_10_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_10_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_10_V_read[21]);
wire tmp_10_22;
assign tmp_10_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_10_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_10_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_10_V_read[22]);
wire tmp_10_23;
assign tmp_10_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_10_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_10_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_10_V_read[23]);
wire tmp_10_24;
assign tmp_10_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_10_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_10_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_10_V_read[24]);
wire tmp_10_25;
assign tmp_10_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_10_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_10_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_10_V_read[25]);
wire tmp_10_26;
assign tmp_10_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_10_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_10_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_10_V_read[26]);
wire tmp_10_27;
assign tmp_10_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_10_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_10_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_10_V_read[27]);
wire tmp_10_28;
assign tmp_10_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_10_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_10_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_10_V_read[28]);
wire tmp_10_29;
assign tmp_10_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_10_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_10_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_10_V_read[29]);
wire tmp_10_30;
assign tmp_10_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_10_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_10_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_10_V_read[30]);
wire tmp_10_31;
assign tmp_10_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_10_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_10_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_10_V_read[31]);
wire tmp_10_32;
assign tmp_10_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_10_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_10_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_10_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_10_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_10_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_10_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_10_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_10_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_10_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_10_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_10_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_10_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_10_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_10_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_10_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_10_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_10_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_10_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_10_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_10_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_10_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_10_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_10_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_10_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_10_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_10_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_10_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_10_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_10_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_10_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_10_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_10_V_read[32]);
wire tmp_10_33;
assign tmp_10_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_10_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_10_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_10_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_10_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_10_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_10_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_10_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_10_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_10_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_10_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_10_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_10_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_10_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_10_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_10_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_10_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_10_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_10_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_10_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_10_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_10_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_10_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_10_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_10_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_10_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_10_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_10_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_10_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_10_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_10_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_10_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_10_V_read[33]);
wire tmp_10_34;
assign tmp_10_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_10_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_10_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_10_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_10_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_10_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_10_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_10_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_10_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_10_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_10_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_10_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_10_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_10_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_10_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_10_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_10_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_10_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_10_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_10_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_10_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_10_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_10_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_10_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_10_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_10_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_10_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_10_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_10_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_10_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_10_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_10_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_10_V_read[34]);
wire tmp_10_35;
assign tmp_10_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_10_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_10_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_10_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_10_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_10_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_10_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_10_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_10_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_10_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_10_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_10_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_10_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_10_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_10_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_10_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_10_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_10_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_10_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_10_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_10_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_10_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_10_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_10_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_10_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_10_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_10_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_10_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_10_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_10_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_10_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_10_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_10_V_read[35]);
wire tmp_10_36;
assign tmp_10_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_10_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_10_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_10_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_10_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_10_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_10_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_10_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_10_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_10_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_10_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_10_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_10_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_10_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_10_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_10_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_10_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_10_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_10_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_10_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_10_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_10_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_10_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_10_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_10_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_10_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_10_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_10_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_10_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_10_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_10_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_10_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_10_V_read[36]);
wire tmp_10_37;
assign tmp_10_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_10_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_10_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_10_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_10_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_10_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_10_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_10_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_10_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_10_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_10_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_10_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_10_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_10_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_10_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_10_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_10_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_10_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_10_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_10_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_10_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_10_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_10_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_10_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_10_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_10_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_10_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_10_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_10_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_10_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_10_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_10_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_10_V_read[37]);
wire tmp_10_38;
assign tmp_10_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_10_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_10_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_10_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_10_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_10_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_10_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_10_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_10_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_10_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_10_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_10_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_10_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_10_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_10_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_10_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_10_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_10_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_10_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_10_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_10_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_10_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_10_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_10_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_10_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_10_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_10_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_10_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_10_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_10_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_10_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_10_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_10_V_read[38]);
wire tmp_10_40;
assign tmp_10_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_10_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_10_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_10_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_10_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_10_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_10_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_10_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_10_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_10_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_10_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_10_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_10_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_10_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_10_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_10_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_10_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_10_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_10_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_10_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_10_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_10_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_10_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_10_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_10_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_10_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_10_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_10_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_10_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_10_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_10_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_10_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_10_V_read[40]);
wire tmp_10_41;
assign tmp_10_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_10_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_10_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_10_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_10_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_10_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_10_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_10_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_10_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_10_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_10_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_10_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_10_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_10_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_10_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_10_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_10_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_10_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_10_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_10_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_10_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_10_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_10_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_10_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_10_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_10_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_10_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_10_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_10_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_10_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_10_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_10_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_10_V_read[41]);
wire tmp_10_42;
assign tmp_10_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_10_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_10_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_10_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_10_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_10_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_10_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_10_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_10_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_10_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_10_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_10_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_10_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_10_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_10_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_10_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_10_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_10_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_10_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_10_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_10_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_10_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_10_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_10_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_10_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_10_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_10_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_10_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_10_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_10_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_10_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_10_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_10_V_read[42]);
wire tmp_10_43;
assign tmp_10_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_10_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_10_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_10_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_10_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_10_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_10_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_10_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_10_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_10_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_10_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_10_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_10_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_10_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_10_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_10_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_10_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_10_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_10_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_10_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_10_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_10_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_10_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_10_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_10_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_10_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_10_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_10_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_10_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_10_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_10_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_10_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_10_V_read[43]);
wire tmp_10_45;
assign tmp_10_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_10_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_10_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_10_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_10_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_10_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_10_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_10_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_10_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_10_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_10_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_10_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_10_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_10_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_10_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_10_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_10_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_10_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_10_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_10_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_10_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_10_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_10_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_10_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_10_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_10_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_10_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_10_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_10_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_10_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_10_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_10_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_10_V_read[45]);
wire tmp_10_47;
assign tmp_10_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_10_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_10_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_10_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_10_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_10_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_10_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_10_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_10_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_10_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_10_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_10_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_10_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_10_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_10_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_10_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_10_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_10_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_10_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_10_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_10_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_10_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_10_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_10_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_10_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_10_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_10_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_10_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_10_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_10_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_10_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_10_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_10_V_read[47]);
wire tmp_10_48;
assign tmp_10_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_10_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_10_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_10_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_10_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_10_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_10_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_10_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_10_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_10_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_10_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_10_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_10_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_10_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_10_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_10_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_10_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_10_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_10_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_10_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_10_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_10_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_10_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_10_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_10_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_10_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_10_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_10_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_10_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_10_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_10_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_10_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_10_V_read[48]);
wire tmp_10_50;
assign tmp_10_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_10_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_10_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_10_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_10_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_10_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_10_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_10_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_10_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_10_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_10_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_10_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_10_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_10_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_10_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_10_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_10_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_10_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_10_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_10_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_10_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_10_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_10_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_10_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_10_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_10_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_10_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_10_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_10_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_10_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_10_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_10_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_10_V_read[50]);
wire tmp_10_51;
assign tmp_10_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_10_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_10_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_10_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_10_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_10_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_10_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_10_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_10_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_10_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_10_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_10_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_10_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_10_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_10_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_10_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_10_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_10_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_10_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_10_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_10_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_10_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_10_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_10_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_10_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_10_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_10_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_10_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_10_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_10_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_10_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_10_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_10_V_read[51]);
wire tmp_10_52;
assign tmp_10_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_10_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_10_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_10_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_10_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_10_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_10_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_10_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_10_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_10_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_10_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_10_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_10_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_10_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_10_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_10_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_10_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_10_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_10_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_10_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_10_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_10_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_10_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_10_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_10_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_10_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_10_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_10_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_10_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_10_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_10_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_10_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_10_V_read[52]);
wire tmp_10_53;
assign tmp_10_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_10_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_10_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_10_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_10_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_10_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_10_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_10_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_10_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_10_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_10_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_10_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_10_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_10_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_10_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_10_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_10_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_10_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_10_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_10_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_10_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_10_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_10_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_10_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_10_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_10_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_10_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_10_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_10_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_10_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_10_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_10_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_10_V_read[53]);
wire tmp_10_56;
assign tmp_10_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_10_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_10_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_10_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_10_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_10_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_10_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_10_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_10_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_10_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_10_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_10_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_10_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_10_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_10_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_10_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_10_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_10_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_10_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_10_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_10_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_10_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_10_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_10_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_10_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_10_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_10_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_10_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_10_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_10_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_10_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_10_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_10_V_read[56]);
wire tmp_10_57;
assign tmp_10_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_10_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_10_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_10_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_10_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_10_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_10_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_10_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_10_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_10_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_10_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_10_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_10_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_10_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_10_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_10_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_10_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_10_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_10_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_10_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_10_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_10_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_10_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_10_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_10_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_10_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_10_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_10_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_10_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_10_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_10_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_10_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_10_V_read[57]);
wire tmp_10_58;
assign tmp_10_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_10_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_10_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_10_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_10_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_10_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_10_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_10_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_10_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_10_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_10_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_10_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_10_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_10_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_10_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_10_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_10_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_10_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_10_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_10_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_10_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_10_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_10_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_10_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_10_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_10_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_10_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_10_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_10_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_10_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_10_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_10_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_10_V_read[58]);
wire tmp_10_59;
assign tmp_10_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_10_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_10_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_10_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_10_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_10_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_10_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_10_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_10_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_10_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_10_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_10_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_10_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_10_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_10_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_10_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_10_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_10_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_10_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_10_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_10_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_10_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_10_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_10_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_10_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_10_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_10_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_10_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_10_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_10_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_10_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_10_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_10_V_read[59]);
wire tmp_10_61;
assign tmp_10_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_10_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_10_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_10_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_10_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_10_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_10_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_10_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_10_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_10_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_10_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_10_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_10_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_10_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_10_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_10_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_10_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_10_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_10_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_10_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_10_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_10_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_10_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_10_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_10_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_10_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_10_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_10_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_10_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_10_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_10_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_10_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_10_V_read[61]);
wire tmp_10_62;
assign tmp_10_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_10_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_10_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_10_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_10_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_10_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_10_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_10_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_10_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_10_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_10_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_10_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_10_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_10_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_10_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_10_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_10_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_10_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_10_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_10_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_10_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_10_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_10_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_10_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_10_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_10_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_10_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_10_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_10_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_10_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_10_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_10_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_10_V_read[62]);
wire tmp_10_64;
assign tmp_10_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_10_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_10_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_10_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_10_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_10_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_10_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_10_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_10_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_10_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_10_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_10_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_10_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_10_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_10_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_10_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_10_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_10_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_10_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_10_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_10_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_10_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_10_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_10_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_10_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_10_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_10_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_10_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_10_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_10_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_10_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_10_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_10_V_read[64]);
wire tmp_10_65;
assign tmp_10_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_10_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_10_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_10_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_10_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_10_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_10_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_10_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_10_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_10_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_10_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_10_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_10_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_10_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_10_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_10_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_10_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_10_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_10_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_10_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_10_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_10_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_10_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_10_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_10_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_10_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_10_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_10_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_10_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_10_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_10_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_10_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_10_V_read[65]);
wire tmp_10_66;
assign tmp_10_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_10_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_10_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_10_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_10_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_10_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_10_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_10_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_10_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_10_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_10_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_10_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_10_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_10_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_10_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_10_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_10_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_10_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_10_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_10_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_10_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_10_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_10_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_10_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_10_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_10_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_10_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_10_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_10_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_10_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_10_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_10_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_10_V_read[66]);
wire tmp_10_67;
assign tmp_10_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_10_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_10_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_10_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_10_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_10_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_10_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_10_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_10_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_10_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_10_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_10_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_10_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_10_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_10_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_10_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_10_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_10_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_10_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_10_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_10_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_10_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_10_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_10_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_10_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_10_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_10_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_10_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_10_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_10_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_10_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_10_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_10_V_read[67]);
wire tmp_10_68;
assign tmp_10_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_10_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_10_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_10_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_10_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_10_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_10_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_10_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_10_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_10_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_10_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_10_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_10_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_10_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_10_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_10_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_10_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_10_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_10_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_10_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_10_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_10_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_10_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_10_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_10_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_10_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_10_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_10_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_10_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_10_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_10_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_10_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_10_V_read[68]);
wire tmp_10_69;
assign tmp_10_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_10_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_10_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_10_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_10_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_10_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_10_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_10_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_10_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_10_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_10_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_10_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_10_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_10_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_10_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_10_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_10_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_10_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_10_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_10_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_10_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_10_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_10_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_10_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_10_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_10_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_10_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_10_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_10_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_10_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_10_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_10_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_10_V_read[69]);
wire tmp_10_70;
assign tmp_10_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_10_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_10_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_10_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_10_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_10_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_10_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_10_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_10_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_10_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_10_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_10_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_10_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_10_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_10_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_10_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_10_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_10_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_10_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_10_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_10_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_10_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_10_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_10_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_10_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_10_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_10_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_10_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_10_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_10_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_10_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_10_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_10_V_read[70]);
wire tmp_10_71;
assign tmp_10_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_10_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_10_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_10_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_10_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_10_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_10_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_10_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_10_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_10_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_10_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_10_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_10_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_10_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_10_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_10_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_10_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_10_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_10_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_10_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_10_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_10_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_10_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_10_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_10_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_10_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_10_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_10_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_10_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_10_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_10_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_10_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_10_V_read[71]);
assign ap_return_10 = {tmp_10_0,tmp_10_1,tmp_10_2,tmp_10_3,tmp_10_4,tmp_10_5,tmp_10_6,tmp_10_7,tmp_10_8,tmp_10_9,tmp_10_10,tmp_10_11,tmp_10_12,tmp_10_13,tmp_10_14,tmp_10_15,tmp_10_16,tmp_10_17,1'b0,tmp_10_19,tmp_10_20,tmp_10_21,tmp_10_22,tmp_10_23,tmp_10_24,tmp_10_25,tmp_10_26,tmp_10_27,tmp_10_28,tmp_10_29,tmp_10_30,tmp_10_31,tmp_10_32,tmp_10_33,tmp_10_34,tmp_10_35,tmp_10_36,tmp_10_37,tmp_10_38,1'b0,tmp_10_40,tmp_10_41,tmp_10_42,tmp_10_43,1'b0,tmp_10_45,1'b0,tmp_10_47,tmp_10_48,1'b0,tmp_10_50,tmp_10_51,tmp_10_52,tmp_10_53,1'b0,1'b0,tmp_10_56,tmp_10_57,tmp_10_58,tmp_10_59,1'b0,tmp_10_61,tmp_10_62,1'b0,tmp_10_64,tmp_10_65,tmp_10_66,tmp_10_67,tmp_10_68,tmp_10_69,tmp_10_70,tmp_10_71};
wire tmp_11_0;
assign tmp_11_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_11_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_11_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_11_V_read[0]);
wire tmp_11_1;
assign tmp_11_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_11_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_11_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_11_V_read[1]);
wire tmp_11_2;
assign tmp_11_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_11_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_11_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_11_V_read[2]);
wire tmp_11_3;
assign tmp_11_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_11_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_11_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_11_V_read[3]);
wire tmp_11_4;
assign tmp_11_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_11_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_11_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_11_V_read[4]);
wire tmp_11_5;
assign tmp_11_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_11_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_11_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_11_V_read[5]);
wire tmp_11_6;
assign tmp_11_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_11_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_11_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_11_V_read[6]);
wire tmp_11_7;
assign tmp_11_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_11_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_11_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_11_V_read[7]);
wire tmp_11_8;
assign tmp_11_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_11_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_11_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_11_V_read[8]);
wire tmp_11_9;
assign tmp_11_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_11_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_11_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_11_V_read[9]);
wire tmp_11_10;
assign tmp_11_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_11_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_11_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_11_V_read[10]);
wire tmp_11_11;
assign tmp_11_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_11_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_11_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_11_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_11_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_11_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_11_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_11_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_11_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_11_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_11_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_11_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_11_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_11_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_11_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_11_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_11_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_11_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_11_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_11_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_11_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_11_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_11_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_11_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_11_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_11_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_11_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_11_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_11_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_11_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_11_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_11_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_11_V_read[11]);
wire tmp_11_12;
assign tmp_11_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_11_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_11_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_11_V_read[12]);
wire tmp_11_13;
assign tmp_11_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_11_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_11_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_11_V_read[13]);
wire tmp_11_14;
assign tmp_11_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_11_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_11_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_11_V_read[14]);
wire tmp_11_15;
assign tmp_11_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_11_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_11_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_11_V_read[15]);
wire tmp_11_16;
assign tmp_11_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_11_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_11_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_11_V_read[16]);
wire tmp_11_17;
assign tmp_11_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_11_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_11_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_11_V_read[17]);
wire tmp_11_18;
assign tmp_11_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_11_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_11_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_11_V_read[18]);
wire tmp_11_19;
assign tmp_11_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_11_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_11_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_11_V_read[19]);
wire tmp_11_20;
assign tmp_11_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_11_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_11_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_11_V_read[20]);
wire tmp_11_21;
assign tmp_11_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_11_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_11_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_11_V_read[21]);
wire tmp_11_22;
assign tmp_11_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_11_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_11_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_11_V_read[22]);
wire tmp_11_24;
assign tmp_11_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_11_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_11_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_11_V_read[24]);
wire tmp_11_26;
assign tmp_11_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_11_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_11_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_11_V_read[26]);
wire tmp_11_27;
assign tmp_11_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_11_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_11_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_11_V_read[27]);
wire tmp_11_28;
assign tmp_11_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_11_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_11_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_11_V_read[28]);
wire tmp_11_29;
assign tmp_11_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_11_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_11_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_11_V_read[29]);
wire tmp_11_30;
assign tmp_11_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_11_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_11_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_11_V_read[30]);
wire tmp_11_31;
assign tmp_11_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_11_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_11_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_11_V_read[31]);
wire tmp_11_32;
assign tmp_11_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_11_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_11_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_11_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_11_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_11_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_11_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_11_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_11_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_11_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_11_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_11_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_11_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_11_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_11_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_11_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_11_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_11_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_11_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_11_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_11_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_11_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_11_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_11_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_11_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_11_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_11_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_11_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_11_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_11_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_11_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_11_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_11_V_read[32]);
wire tmp_11_33;
assign tmp_11_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_11_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_11_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_11_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_11_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_11_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_11_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_11_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_11_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_11_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_11_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_11_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_11_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_11_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_11_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_11_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_11_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_11_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_11_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_11_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_11_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_11_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_11_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_11_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_11_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_11_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_11_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_11_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_11_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_11_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_11_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_11_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_11_V_read[33]);
wire tmp_11_34;
assign tmp_11_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_11_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_11_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_11_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_11_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_11_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_11_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_11_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_11_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_11_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_11_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_11_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_11_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_11_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_11_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_11_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_11_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_11_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_11_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_11_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_11_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_11_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_11_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_11_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_11_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_11_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_11_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_11_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_11_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_11_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_11_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_11_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_11_V_read[34]);
wire tmp_11_35;
assign tmp_11_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_11_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_11_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_11_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_11_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_11_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_11_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_11_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_11_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_11_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_11_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_11_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_11_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_11_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_11_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_11_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_11_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_11_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_11_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_11_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_11_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_11_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_11_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_11_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_11_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_11_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_11_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_11_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_11_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_11_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_11_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_11_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_11_V_read[35]);
wire tmp_11_36;
assign tmp_11_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_11_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_11_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_11_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_11_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_11_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_11_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_11_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_11_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_11_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_11_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_11_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_11_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_11_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_11_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_11_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_11_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_11_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_11_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_11_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_11_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_11_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_11_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_11_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_11_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_11_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_11_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_11_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_11_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_11_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_11_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_11_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_11_V_read[36]);
wire tmp_11_37;
assign tmp_11_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_11_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_11_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_11_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_11_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_11_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_11_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_11_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_11_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_11_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_11_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_11_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_11_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_11_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_11_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_11_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_11_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_11_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_11_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_11_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_11_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_11_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_11_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_11_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_11_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_11_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_11_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_11_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_11_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_11_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_11_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_11_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_11_V_read[37]);
wire tmp_11_38;
assign tmp_11_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_11_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_11_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_11_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_11_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_11_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_11_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_11_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_11_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_11_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_11_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_11_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_11_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_11_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_11_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_11_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_11_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_11_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_11_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_11_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_11_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_11_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_11_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_11_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_11_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_11_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_11_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_11_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_11_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_11_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_11_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_11_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_11_V_read[38]);
wire tmp_11_40;
assign tmp_11_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_11_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_11_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_11_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_11_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_11_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_11_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_11_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_11_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_11_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_11_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_11_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_11_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_11_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_11_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_11_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_11_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_11_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_11_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_11_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_11_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_11_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_11_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_11_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_11_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_11_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_11_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_11_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_11_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_11_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_11_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_11_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_11_V_read[40]);
wire tmp_11_41;
assign tmp_11_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_11_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_11_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_11_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_11_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_11_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_11_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_11_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_11_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_11_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_11_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_11_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_11_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_11_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_11_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_11_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_11_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_11_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_11_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_11_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_11_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_11_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_11_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_11_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_11_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_11_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_11_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_11_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_11_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_11_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_11_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_11_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_11_V_read[41]);
wire tmp_11_42;
assign tmp_11_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_11_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_11_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_11_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_11_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_11_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_11_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_11_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_11_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_11_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_11_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_11_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_11_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_11_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_11_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_11_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_11_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_11_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_11_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_11_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_11_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_11_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_11_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_11_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_11_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_11_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_11_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_11_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_11_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_11_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_11_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_11_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_11_V_read[42]);
wire tmp_11_43;
assign tmp_11_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_11_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_11_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_11_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_11_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_11_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_11_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_11_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_11_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_11_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_11_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_11_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_11_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_11_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_11_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_11_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_11_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_11_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_11_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_11_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_11_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_11_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_11_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_11_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_11_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_11_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_11_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_11_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_11_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_11_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_11_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_11_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_11_V_read[43]);
wire tmp_11_44;
assign tmp_11_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_11_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_11_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_11_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_11_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_11_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_11_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_11_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_11_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_11_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_11_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_11_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_11_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_11_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_11_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_11_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_11_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_11_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_11_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_11_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_11_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_11_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_11_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_11_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_11_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_11_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_11_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_11_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_11_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_11_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_11_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_11_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_11_V_read[44]);
wire tmp_11_45;
assign tmp_11_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_11_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_11_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_11_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_11_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_11_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_11_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_11_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_11_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_11_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_11_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_11_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_11_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_11_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_11_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_11_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_11_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_11_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_11_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_11_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_11_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_11_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_11_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_11_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_11_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_11_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_11_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_11_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_11_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_11_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_11_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_11_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_11_V_read[45]);
wire tmp_11_46;
assign tmp_11_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_11_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_11_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_11_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_11_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_11_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_11_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_11_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_11_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_11_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_11_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_11_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_11_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_11_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_11_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_11_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_11_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_11_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_11_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_11_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_11_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_11_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_11_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_11_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_11_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_11_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_11_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_11_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_11_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_11_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_11_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_11_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_11_V_read[46]);
wire tmp_11_48;
assign tmp_11_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_11_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_11_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_11_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_11_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_11_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_11_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_11_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_11_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_11_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_11_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_11_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_11_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_11_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_11_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_11_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_11_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_11_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_11_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_11_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_11_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_11_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_11_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_11_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_11_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_11_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_11_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_11_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_11_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_11_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_11_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_11_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_11_V_read[48]);
wire tmp_11_49;
assign tmp_11_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_11_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_11_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_11_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_11_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_11_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_11_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_11_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_11_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_11_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_11_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_11_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_11_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_11_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_11_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_11_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_11_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_11_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_11_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_11_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_11_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_11_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_11_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_11_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_11_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_11_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_11_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_11_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_11_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_11_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_11_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_11_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_11_V_read[49]);
wire tmp_11_50;
assign tmp_11_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_11_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_11_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_11_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_11_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_11_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_11_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_11_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_11_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_11_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_11_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_11_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_11_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_11_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_11_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_11_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_11_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_11_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_11_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_11_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_11_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_11_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_11_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_11_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_11_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_11_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_11_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_11_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_11_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_11_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_11_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_11_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_11_V_read[50]);
wire tmp_11_51;
assign tmp_11_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_11_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_11_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_11_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_11_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_11_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_11_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_11_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_11_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_11_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_11_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_11_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_11_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_11_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_11_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_11_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_11_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_11_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_11_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_11_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_11_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_11_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_11_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_11_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_11_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_11_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_11_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_11_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_11_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_11_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_11_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_11_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_11_V_read[51]);
wire tmp_11_52;
assign tmp_11_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_11_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_11_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_11_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_11_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_11_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_11_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_11_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_11_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_11_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_11_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_11_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_11_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_11_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_11_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_11_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_11_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_11_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_11_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_11_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_11_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_11_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_11_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_11_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_11_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_11_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_11_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_11_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_11_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_11_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_11_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_11_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_11_V_read[52]);
wire tmp_11_54;
assign tmp_11_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_11_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_11_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_11_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_11_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_11_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_11_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_11_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_11_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_11_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_11_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_11_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_11_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_11_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_11_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_11_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_11_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_11_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_11_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_11_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_11_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_11_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_11_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_11_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_11_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_11_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_11_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_11_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_11_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_11_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_11_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_11_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_11_V_read[54]);
wire tmp_11_55;
assign tmp_11_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_11_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_11_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_11_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_11_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_11_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_11_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_11_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_11_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_11_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_11_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_11_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_11_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_11_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_11_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_11_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_11_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_11_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_11_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_11_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_11_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_11_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_11_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_11_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_11_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_11_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_11_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_11_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_11_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_11_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_11_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_11_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_11_V_read[55]);
wire tmp_11_56;
assign tmp_11_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_11_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_11_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_11_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_11_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_11_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_11_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_11_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_11_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_11_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_11_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_11_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_11_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_11_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_11_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_11_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_11_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_11_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_11_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_11_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_11_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_11_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_11_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_11_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_11_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_11_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_11_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_11_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_11_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_11_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_11_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_11_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_11_V_read[56]);
wire tmp_11_57;
assign tmp_11_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_11_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_11_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_11_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_11_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_11_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_11_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_11_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_11_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_11_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_11_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_11_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_11_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_11_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_11_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_11_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_11_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_11_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_11_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_11_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_11_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_11_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_11_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_11_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_11_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_11_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_11_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_11_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_11_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_11_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_11_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_11_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_11_V_read[57]);
wire tmp_11_59;
assign tmp_11_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_11_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_11_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_11_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_11_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_11_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_11_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_11_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_11_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_11_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_11_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_11_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_11_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_11_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_11_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_11_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_11_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_11_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_11_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_11_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_11_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_11_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_11_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_11_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_11_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_11_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_11_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_11_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_11_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_11_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_11_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_11_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_11_V_read[59]);
wire tmp_11_60;
assign tmp_11_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_11_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_11_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_11_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_11_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_11_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_11_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_11_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_11_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_11_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_11_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_11_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_11_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_11_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_11_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_11_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_11_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_11_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_11_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_11_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_11_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_11_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_11_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_11_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_11_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_11_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_11_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_11_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_11_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_11_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_11_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_11_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_11_V_read[60]);
wire tmp_11_61;
assign tmp_11_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_11_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_11_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_11_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_11_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_11_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_11_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_11_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_11_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_11_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_11_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_11_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_11_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_11_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_11_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_11_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_11_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_11_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_11_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_11_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_11_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_11_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_11_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_11_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_11_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_11_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_11_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_11_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_11_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_11_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_11_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_11_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_11_V_read[61]);
wire tmp_11_62;
assign tmp_11_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_11_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_11_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_11_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_11_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_11_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_11_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_11_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_11_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_11_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_11_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_11_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_11_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_11_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_11_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_11_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_11_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_11_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_11_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_11_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_11_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_11_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_11_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_11_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_11_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_11_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_11_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_11_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_11_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_11_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_11_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_11_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_11_V_read[62]);
wire tmp_11_63;
assign tmp_11_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_11_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_11_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_11_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_11_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_11_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_11_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_11_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_11_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_11_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_11_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_11_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_11_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_11_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_11_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_11_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_11_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_11_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_11_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_11_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_11_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_11_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_11_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_11_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_11_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_11_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_11_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_11_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_11_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_11_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_11_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_11_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_11_V_read[63]);
wire tmp_11_64;
assign tmp_11_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_11_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_11_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_11_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_11_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_11_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_11_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_11_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_11_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_11_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_11_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_11_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_11_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_11_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_11_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_11_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_11_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_11_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_11_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_11_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_11_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_11_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_11_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_11_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_11_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_11_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_11_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_11_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_11_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_11_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_11_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_11_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_11_V_read[64]);
wire tmp_11_65;
assign tmp_11_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_11_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_11_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_11_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_11_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_11_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_11_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_11_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_11_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_11_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_11_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_11_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_11_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_11_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_11_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_11_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_11_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_11_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_11_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_11_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_11_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_11_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_11_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_11_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_11_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_11_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_11_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_11_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_11_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_11_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_11_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_11_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_11_V_read[65]);
wire tmp_11_66;
assign tmp_11_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_11_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_11_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_11_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_11_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_11_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_11_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_11_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_11_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_11_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_11_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_11_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_11_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_11_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_11_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_11_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_11_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_11_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_11_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_11_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_11_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_11_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_11_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_11_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_11_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_11_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_11_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_11_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_11_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_11_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_11_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_11_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_11_V_read[66]);
wire tmp_11_67;
assign tmp_11_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_11_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_11_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_11_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_11_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_11_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_11_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_11_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_11_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_11_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_11_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_11_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_11_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_11_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_11_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_11_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_11_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_11_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_11_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_11_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_11_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_11_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_11_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_11_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_11_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_11_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_11_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_11_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_11_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_11_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_11_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_11_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_11_V_read[67]);
wire tmp_11_68;
assign tmp_11_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_11_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_11_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_11_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_11_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_11_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_11_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_11_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_11_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_11_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_11_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_11_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_11_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_11_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_11_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_11_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_11_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_11_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_11_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_11_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_11_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_11_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_11_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_11_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_11_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_11_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_11_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_11_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_11_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_11_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_11_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_11_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_11_V_read[68]);
wire tmp_11_69;
assign tmp_11_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_11_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_11_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_11_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_11_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_11_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_11_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_11_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_11_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_11_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_11_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_11_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_11_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_11_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_11_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_11_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_11_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_11_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_11_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_11_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_11_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_11_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_11_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_11_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_11_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_11_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_11_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_11_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_11_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_11_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_11_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_11_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_11_V_read[69]);
wire tmp_11_70;
assign tmp_11_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_11_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_11_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_11_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_11_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_11_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_11_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_11_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_11_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_11_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_11_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_11_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_11_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_11_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_11_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_11_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_11_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_11_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_11_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_11_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_11_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_11_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_11_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_11_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_11_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_11_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_11_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_11_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_11_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_11_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_11_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_11_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_11_V_read[70]);
assign ap_return_11 = {tmp_11_0,tmp_11_1,tmp_11_2,tmp_11_3,tmp_11_4,tmp_11_5,tmp_11_6,tmp_11_7,tmp_11_8,tmp_11_9,tmp_11_10,tmp_11_11,tmp_11_12,tmp_11_13,tmp_11_14,tmp_11_15,tmp_11_16,tmp_11_17,tmp_11_18,tmp_11_19,tmp_11_20,tmp_11_21,tmp_11_22,1'b0,tmp_11_24,1'b0,tmp_11_26,tmp_11_27,tmp_11_28,tmp_11_29,tmp_11_30,tmp_11_31,tmp_11_32,tmp_11_33,tmp_11_34,tmp_11_35,tmp_11_36,tmp_11_37,tmp_11_38,1'b0,tmp_11_40,tmp_11_41,tmp_11_42,tmp_11_43,tmp_11_44,tmp_11_45,tmp_11_46,1'b0,tmp_11_48,tmp_11_49,tmp_11_50,tmp_11_51,tmp_11_52,1'b0,tmp_11_54,tmp_11_55,tmp_11_56,tmp_11_57,1'b0,tmp_11_59,tmp_11_60,tmp_11_61,tmp_11_62,tmp_11_63,tmp_11_64,tmp_11_65,tmp_11_66,tmp_11_67,tmp_11_68,tmp_11_69,tmp_11_70,1'b0};
wire tmp_12_0;
assign tmp_12_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_12_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_12_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_12_V_read[0]);
wire tmp_12_1;
assign tmp_12_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_12_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_12_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_12_V_read[1]);
wire tmp_12_2;
assign tmp_12_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_12_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_12_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_12_V_read[2]);
wire tmp_12_3;
assign tmp_12_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_12_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_12_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_12_V_read[3]);
wire tmp_12_4;
assign tmp_12_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_12_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_12_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_12_V_read[4]);
wire tmp_12_5;
assign tmp_12_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_12_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_12_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_12_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_12_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_12_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_12_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_12_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_12_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_12_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_12_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_12_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_12_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_12_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_12_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_12_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_12_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_12_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_12_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_12_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_12_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_12_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_12_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_12_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_12_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_12_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_12_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_12_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_12_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_12_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_12_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_12_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_12_V_read[5]);
wire tmp_12_6;
assign tmp_12_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_12_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_12_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_12_V_read[6]);
wire tmp_12_7;
assign tmp_12_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_12_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_12_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_12_V_read[7]);
wire tmp_12_8;
assign tmp_12_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_12_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_12_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_12_V_read[8]);
wire tmp_12_9;
assign tmp_12_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_12_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_12_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_12_V_read[9]);
wire tmp_12_10;
assign tmp_12_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_12_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_12_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_12_V_read[10]);
wire tmp_12_11;
assign tmp_12_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_12_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_12_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_12_V_read[11]);
wire tmp_12_12;
assign tmp_12_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_12_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_12_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_12_V_read[12]);
wire tmp_12_13;
assign tmp_12_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_12_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_12_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_12_V_read[13]);
wire tmp_12_14;
assign tmp_12_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_12_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_12_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_12_V_read[14]);
wire tmp_12_15;
assign tmp_12_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_12_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_12_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_12_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_12_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_12_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_12_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_12_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_12_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_12_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_12_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_12_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_12_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_12_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_12_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_12_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_12_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_12_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_12_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_12_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_12_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_12_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_12_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_12_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_12_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_12_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_12_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_12_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_12_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_12_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_12_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_12_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_12_V_read[15]);
wire tmp_12_16;
assign tmp_12_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_12_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_12_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_12_V_read[16]);
wire tmp_12_17;
assign tmp_12_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_12_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_12_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_12_V_read[17]);
wire tmp_12_18;
assign tmp_12_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_12_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_12_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_12_V_read[18]);
wire tmp_12_19;
assign tmp_12_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_12_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_12_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_12_V_read[19]);
wire tmp_12_20;
assign tmp_12_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_12_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_12_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_12_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_12_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_12_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_12_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_12_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_12_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_12_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_12_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_12_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_12_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_12_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_12_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_12_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_12_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_12_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_12_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_12_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_12_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_12_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_12_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_12_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_12_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_12_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_12_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_12_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_12_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_12_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_12_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_12_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_12_V_read[20]);
wire tmp_12_21;
assign tmp_12_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_12_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_12_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_12_V_read[21]);
wire tmp_12_22;
assign tmp_12_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_12_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_12_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_12_V_read[22]);
wire tmp_12_23;
assign tmp_12_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_12_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_12_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_12_V_read[23]);
wire tmp_12_24;
assign tmp_12_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_12_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_12_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_12_V_read[24]);
wire tmp_12_25;
assign tmp_12_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_12_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_12_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_12_V_read[25]);
wire tmp_12_26;
assign tmp_12_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_12_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_12_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_12_V_read[26]);
wire tmp_12_27;
assign tmp_12_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_12_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_12_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_12_V_read[27]);
wire tmp_12_28;
assign tmp_12_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_12_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_12_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_12_V_read[28]);
wire tmp_12_29;
assign tmp_12_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_12_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_12_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_12_V_read[29]);
wire tmp_12_30;
assign tmp_12_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_12_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_12_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_12_V_read[30]);
wire tmp_12_31;
assign tmp_12_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_12_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_12_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_12_V_read[31]);
wire tmp_12_32;
assign tmp_12_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_12_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_12_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_12_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_12_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_12_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_12_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_12_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_12_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_12_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_12_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_12_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_12_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_12_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_12_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_12_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_12_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_12_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_12_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_12_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_12_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_12_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_12_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_12_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_12_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_12_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_12_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_12_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_12_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_12_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_12_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_12_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_12_V_read[32]);
wire tmp_12_33;
assign tmp_12_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_12_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_12_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_12_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_12_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_12_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_12_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_12_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_12_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_12_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_12_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_12_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_12_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_12_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_12_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_12_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_12_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_12_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_12_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_12_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_12_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_12_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_12_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_12_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_12_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_12_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_12_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_12_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_12_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_12_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_12_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_12_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_12_V_read[33]);
wire tmp_12_34;
assign tmp_12_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_12_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_12_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_12_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_12_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_12_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_12_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_12_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_12_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_12_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_12_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_12_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_12_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_12_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_12_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_12_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_12_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_12_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_12_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_12_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_12_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_12_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_12_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_12_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_12_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_12_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_12_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_12_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_12_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_12_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_12_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_12_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_12_V_read[34]);
wire tmp_12_35;
assign tmp_12_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_12_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_12_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_12_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_12_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_12_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_12_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_12_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_12_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_12_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_12_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_12_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_12_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_12_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_12_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_12_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_12_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_12_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_12_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_12_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_12_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_12_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_12_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_12_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_12_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_12_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_12_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_12_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_12_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_12_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_12_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_12_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_12_V_read[35]);
wire tmp_12_36;
assign tmp_12_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_12_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_12_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_12_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_12_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_12_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_12_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_12_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_12_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_12_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_12_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_12_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_12_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_12_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_12_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_12_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_12_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_12_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_12_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_12_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_12_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_12_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_12_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_12_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_12_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_12_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_12_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_12_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_12_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_12_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_12_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_12_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_12_V_read[36]);
wire tmp_12_38;
assign tmp_12_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_12_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_12_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_12_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_12_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_12_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_12_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_12_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_12_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_12_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_12_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_12_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_12_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_12_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_12_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_12_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_12_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_12_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_12_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_12_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_12_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_12_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_12_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_12_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_12_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_12_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_12_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_12_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_12_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_12_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_12_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_12_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_12_V_read[38]);
wire tmp_12_40;
assign tmp_12_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_12_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_12_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_12_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_12_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_12_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_12_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_12_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_12_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_12_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_12_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_12_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_12_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_12_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_12_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_12_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_12_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_12_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_12_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_12_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_12_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_12_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_12_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_12_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_12_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_12_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_12_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_12_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_12_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_12_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_12_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_12_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_12_V_read[40]);
wire tmp_12_41;
assign tmp_12_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_12_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_12_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_12_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_12_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_12_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_12_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_12_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_12_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_12_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_12_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_12_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_12_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_12_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_12_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_12_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_12_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_12_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_12_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_12_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_12_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_12_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_12_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_12_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_12_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_12_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_12_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_12_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_12_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_12_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_12_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_12_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_12_V_read[41]);
wire tmp_12_42;
assign tmp_12_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_12_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_12_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_12_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_12_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_12_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_12_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_12_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_12_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_12_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_12_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_12_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_12_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_12_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_12_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_12_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_12_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_12_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_12_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_12_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_12_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_12_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_12_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_12_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_12_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_12_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_12_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_12_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_12_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_12_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_12_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_12_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_12_V_read[42]);
wire tmp_12_43;
assign tmp_12_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_12_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_12_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_12_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_12_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_12_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_12_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_12_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_12_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_12_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_12_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_12_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_12_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_12_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_12_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_12_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_12_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_12_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_12_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_12_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_12_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_12_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_12_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_12_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_12_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_12_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_12_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_12_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_12_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_12_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_12_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_12_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_12_V_read[43]);
wire tmp_12_44;
assign tmp_12_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_12_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_12_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_12_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_12_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_12_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_12_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_12_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_12_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_12_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_12_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_12_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_12_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_12_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_12_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_12_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_12_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_12_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_12_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_12_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_12_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_12_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_12_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_12_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_12_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_12_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_12_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_12_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_12_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_12_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_12_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_12_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_12_V_read[44]);
wire tmp_12_45;
assign tmp_12_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_12_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_12_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_12_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_12_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_12_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_12_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_12_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_12_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_12_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_12_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_12_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_12_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_12_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_12_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_12_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_12_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_12_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_12_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_12_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_12_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_12_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_12_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_12_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_12_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_12_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_12_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_12_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_12_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_12_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_12_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_12_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_12_V_read[45]);
wire tmp_12_46;
assign tmp_12_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_12_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_12_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_12_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_12_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_12_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_12_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_12_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_12_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_12_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_12_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_12_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_12_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_12_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_12_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_12_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_12_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_12_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_12_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_12_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_12_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_12_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_12_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_12_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_12_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_12_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_12_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_12_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_12_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_12_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_12_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_12_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_12_V_read[46]);
wire tmp_12_48;
assign tmp_12_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_12_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_12_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_12_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_12_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_12_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_12_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_12_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_12_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_12_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_12_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_12_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_12_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_12_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_12_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_12_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_12_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_12_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_12_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_12_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_12_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_12_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_12_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_12_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_12_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_12_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_12_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_12_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_12_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_12_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_12_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_12_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_12_V_read[48]);
wire tmp_12_49;
assign tmp_12_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_12_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_12_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_12_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_12_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_12_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_12_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_12_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_12_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_12_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_12_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_12_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_12_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_12_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_12_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_12_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_12_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_12_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_12_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_12_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_12_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_12_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_12_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_12_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_12_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_12_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_12_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_12_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_12_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_12_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_12_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_12_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_12_V_read[49]);
wire tmp_12_50;
assign tmp_12_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_12_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_12_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_12_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_12_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_12_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_12_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_12_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_12_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_12_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_12_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_12_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_12_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_12_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_12_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_12_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_12_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_12_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_12_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_12_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_12_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_12_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_12_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_12_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_12_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_12_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_12_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_12_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_12_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_12_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_12_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_12_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_12_V_read[50]);
wire tmp_12_51;
assign tmp_12_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_12_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_12_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_12_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_12_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_12_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_12_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_12_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_12_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_12_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_12_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_12_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_12_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_12_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_12_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_12_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_12_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_12_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_12_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_12_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_12_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_12_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_12_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_12_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_12_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_12_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_12_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_12_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_12_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_12_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_12_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_12_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_12_V_read[51]);
wire tmp_12_53;
assign tmp_12_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_12_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_12_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_12_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_12_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_12_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_12_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_12_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_12_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_12_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_12_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_12_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_12_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_12_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_12_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_12_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_12_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_12_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_12_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_12_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_12_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_12_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_12_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_12_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_12_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_12_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_12_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_12_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_12_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_12_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_12_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_12_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_12_V_read[53]);
wire tmp_12_54;
assign tmp_12_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_12_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_12_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_12_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_12_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_12_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_12_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_12_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_12_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_12_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_12_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_12_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_12_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_12_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_12_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_12_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_12_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_12_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_12_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_12_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_12_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_12_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_12_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_12_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_12_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_12_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_12_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_12_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_12_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_12_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_12_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_12_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_12_V_read[54]);
wire tmp_12_55;
assign tmp_12_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_12_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_12_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_12_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_12_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_12_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_12_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_12_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_12_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_12_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_12_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_12_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_12_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_12_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_12_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_12_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_12_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_12_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_12_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_12_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_12_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_12_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_12_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_12_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_12_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_12_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_12_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_12_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_12_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_12_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_12_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_12_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_12_V_read[55]);
wire tmp_12_56;
assign tmp_12_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_12_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_12_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_12_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_12_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_12_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_12_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_12_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_12_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_12_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_12_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_12_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_12_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_12_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_12_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_12_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_12_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_12_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_12_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_12_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_12_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_12_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_12_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_12_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_12_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_12_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_12_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_12_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_12_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_12_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_12_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_12_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_12_V_read[56]);
wire tmp_12_57;
assign tmp_12_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_12_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_12_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_12_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_12_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_12_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_12_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_12_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_12_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_12_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_12_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_12_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_12_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_12_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_12_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_12_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_12_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_12_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_12_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_12_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_12_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_12_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_12_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_12_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_12_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_12_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_12_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_12_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_12_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_12_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_12_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_12_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_12_V_read[57]);
wire tmp_12_58;
assign tmp_12_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_12_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_12_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_12_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_12_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_12_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_12_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_12_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_12_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_12_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_12_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_12_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_12_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_12_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_12_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_12_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_12_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_12_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_12_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_12_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_12_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_12_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_12_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_12_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_12_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_12_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_12_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_12_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_12_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_12_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_12_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_12_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_12_V_read[58]);
wire tmp_12_60;
assign tmp_12_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_12_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_12_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_12_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_12_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_12_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_12_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_12_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_12_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_12_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_12_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_12_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_12_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_12_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_12_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_12_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_12_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_12_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_12_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_12_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_12_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_12_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_12_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_12_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_12_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_12_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_12_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_12_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_12_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_12_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_12_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_12_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_12_V_read[60]);
wire tmp_12_61;
assign tmp_12_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_12_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_12_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_12_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_12_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_12_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_12_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_12_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_12_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_12_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_12_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_12_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_12_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_12_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_12_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_12_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_12_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_12_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_12_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_12_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_12_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_12_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_12_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_12_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_12_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_12_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_12_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_12_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_12_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_12_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_12_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_12_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_12_V_read[61]);
wire tmp_12_62;
assign tmp_12_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_12_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_12_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_12_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_12_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_12_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_12_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_12_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_12_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_12_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_12_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_12_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_12_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_12_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_12_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_12_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_12_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_12_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_12_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_12_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_12_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_12_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_12_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_12_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_12_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_12_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_12_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_12_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_12_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_12_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_12_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_12_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_12_V_read[62]);
wire tmp_12_63;
assign tmp_12_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_12_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_12_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_12_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_12_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_12_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_12_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_12_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_12_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_12_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_12_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_12_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_12_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_12_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_12_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_12_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_12_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_12_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_12_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_12_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_12_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_12_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_12_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_12_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_12_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_12_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_12_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_12_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_12_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_12_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_12_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_12_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_12_V_read[63]);
wire tmp_12_64;
assign tmp_12_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_12_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_12_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_12_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_12_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_12_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_12_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_12_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_12_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_12_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_12_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_12_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_12_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_12_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_12_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_12_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_12_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_12_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_12_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_12_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_12_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_12_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_12_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_12_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_12_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_12_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_12_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_12_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_12_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_12_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_12_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_12_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_12_V_read[64]);
wire tmp_12_65;
assign tmp_12_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_12_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_12_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_12_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_12_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_12_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_12_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_12_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_12_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_12_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_12_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_12_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_12_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_12_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_12_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_12_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_12_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_12_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_12_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_12_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_12_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_12_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_12_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_12_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_12_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_12_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_12_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_12_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_12_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_12_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_12_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_12_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_12_V_read[65]);
wire tmp_12_66;
assign tmp_12_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_12_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_12_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_12_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_12_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_12_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_12_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_12_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_12_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_12_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_12_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_12_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_12_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_12_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_12_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_12_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_12_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_12_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_12_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_12_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_12_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_12_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_12_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_12_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_12_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_12_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_12_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_12_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_12_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_12_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_12_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_12_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_12_V_read[66]);
wire tmp_12_67;
assign tmp_12_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_12_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_12_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_12_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_12_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_12_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_12_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_12_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_12_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_12_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_12_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_12_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_12_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_12_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_12_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_12_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_12_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_12_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_12_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_12_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_12_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_12_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_12_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_12_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_12_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_12_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_12_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_12_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_12_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_12_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_12_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_12_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_12_V_read[67]);
wire tmp_12_68;
assign tmp_12_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_12_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_12_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_12_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_12_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_12_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_12_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_12_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_12_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_12_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_12_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_12_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_12_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_12_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_12_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_12_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_12_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_12_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_12_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_12_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_12_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_12_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_12_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_12_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_12_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_12_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_12_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_12_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_12_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_12_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_12_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_12_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_12_V_read[68]);
wire tmp_12_69;
assign tmp_12_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_12_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_12_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_12_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_12_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_12_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_12_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_12_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_12_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_12_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_12_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_12_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_12_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_12_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_12_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_12_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_12_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_12_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_12_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_12_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_12_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_12_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_12_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_12_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_12_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_12_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_12_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_12_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_12_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_12_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_12_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_12_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_12_V_read[69]);
wire tmp_12_70;
assign tmp_12_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_12_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_12_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_12_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_12_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_12_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_12_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_12_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_12_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_12_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_12_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_12_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_12_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_12_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_12_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_12_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_12_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_12_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_12_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_12_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_12_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_12_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_12_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_12_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_12_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_12_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_12_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_12_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_12_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_12_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_12_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_12_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_12_V_read[70]);
wire tmp_12_71;
assign tmp_12_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_12_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_12_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_12_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_12_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_12_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_12_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_12_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_12_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_12_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_12_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_12_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_12_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_12_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_12_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_12_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_12_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_12_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_12_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_12_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_12_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_12_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_12_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_12_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_12_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_12_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_12_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_12_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_12_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_12_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_12_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_12_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_12_V_read[71]);
assign ap_return_12 = {tmp_12_0,tmp_12_1,tmp_12_2,tmp_12_3,tmp_12_4,tmp_12_5,tmp_12_6,tmp_12_7,tmp_12_8,tmp_12_9,tmp_12_10,tmp_12_11,tmp_12_12,tmp_12_13,tmp_12_14,tmp_12_15,tmp_12_16,tmp_12_17,tmp_12_18,tmp_12_19,tmp_12_20,tmp_12_21,tmp_12_22,tmp_12_23,tmp_12_24,tmp_12_25,tmp_12_26,tmp_12_27,tmp_12_28,tmp_12_29,tmp_12_30,tmp_12_31,tmp_12_32,tmp_12_33,tmp_12_34,tmp_12_35,tmp_12_36,1'b0,tmp_12_38,1'b0,tmp_12_40,tmp_12_41,tmp_12_42,tmp_12_43,tmp_12_44,tmp_12_45,tmp_12_46,1'b0,tmp_12_48,tmp_12_49,tmp_12_50,tmp_12_51,1'b0,tmp_12_53,tmp_12_54,tmp_12_55,tmp_12_56,tmp_12_57,tmp_12_58,1'b0,tmp_12_60,tmp_12_61,tmp_12_62,tmp_12_63,tmp_12_64,tmp_12_65,tmp_12_66,tmp_12_67,tmp_12_68,tmp_12_69,tmp_12_70,tmp_12_71};
wire tmp_13_0;
assign tmp_13_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_13_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_13_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_13_V_read[0]);
wire tmp_13_1;
assign tmp_13_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_13_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_13_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_13_V_read[1]);
wire tmp_13_2;
assign tmp_13_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_13_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_13_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_13_V_read[2]);
wire tmp_13_3;
assign tmp_13_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_13_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_13_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_13_V_read[3]);
wire tmp_13_4;
assign tmp_13_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_13_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_13_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_13_V_read[4]);
wire tmp_13_5;
assign tmp_13_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_13_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_13_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_13_V_read[5]);
wire tmp_13_7;
assign tmp_13_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_13_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_13_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_13_V_read[7]);
wire tmp_13_8;
assign tmp_13_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_13_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_13_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_13_V_read[8]);
wire tmp_13_9;
assign tmp_13_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_13_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_13_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_13_V_read[9]);
wire tmp_13_10;
assign tmp_13_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_13_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_13_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_13_V_read[10]);
wire tmp_13_11;
assign tmp_13_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_13_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_13_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_13_V_read[11]);
wire tmp_13_12;
assign tmp_13_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_13_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_13_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_13_V_read[12]);
wire tmp_13_13;
assign tmp_13_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_13_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_13_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_13_V_read[13]);
wire tmp_13_14;
assign tmp_13_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_13_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_13_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_13_V_read[14]);
wire tmp_13_15;
assign tmp_13_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_13_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_13_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_13_V_read[15]);
wire tmp_13_16;
assign tmp_13_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_13_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_13_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_13_V_read[16]);
wire tmp_13_17;
assign tmp_13_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_13_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_13_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_13_V_read[17]);
wire tmp_13_18;
assign tmp_13_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_13_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_13_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_13_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_13_V_read[18]);
wire tmp_13_19;
assign tmp_13_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_13_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_13_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_13_V_read[19]);
wire tmp_13_20;
assign tmp_13_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_13_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_13_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_13_V_read[20]);
wire tmp_13_21;
assign tmp_13_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_13_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_13_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_13_V_read[21]);
wire tmp_13_22;
assign tmp_13_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_13_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_13_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_13_V_read[22]);
wire tmp_13_23;
assign tmp_13_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_13_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_13_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_13_V_read[23]);
wire tmp_13_24;
assign tmp_13_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_13_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_13_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_13_V_read[24]);
wire tmp_13_25;
assign tmp_13_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_13_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_13_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_13_V_read[25]);
wire tmp_13_26;
assign tmp_13_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_13_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_13_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_13_V_read[26]);
wire tmp_13_27;
assign tmp_13_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_13_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_13_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_13_V_read[27]);
wire tmp_13_28;
assign tmp_13_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_13_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_13_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_13_V_read[28]);
wire tmp_13_29;
assign tmp_13_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_13_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_13_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_13_V_read[29]);
wire tmp_13_30;
assign tmp_13_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_13_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_13_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_13_V_read[30]);
wire tmp_13_31;
assign tmp_13_31 = (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (1 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (0 &  in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] &  in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] &  in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] &  in_3_V[31] & ~weight_0_13_V_read[31]) | (0 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] &  weight_0_13_V_read[31]) | (1 & ~in_V[31] & ~in_1_V[31] & ~in_2_V[31] & ~in_3_V[31] & ~weight_0_13_V_read[31]);
wire tmp_13_32;
assign tmp_13_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_13_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_13_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_13_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_13_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_13_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_13_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_13_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_13_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_13_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_13_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_13_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_13_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_13_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_13_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_13_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_13_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_13_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_13_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_13_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_13_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_13_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_13_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_13_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_13_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_13_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_13_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_13_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_13_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_13_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_13_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_13_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_13_V_read[32]);
wire tmp_13_33;
assign tmp_13_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_13_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_13_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_13_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_13_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_13_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_13_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_13_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_13_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_13_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_13_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_13_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_13_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_13_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_13_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_13_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_13_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_13_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_13_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_13_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_13_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_13_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_13_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_13_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_13_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_13_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_13_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_13_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_13_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_13_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_13_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_13_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_13_V_read[33]);
wire tmp_13_35;
assign tmp_13_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_13_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_13_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_13_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_13_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_13_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_13_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_13_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_13_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_13_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_13_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_13_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_13_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_13_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_13_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_13_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_13_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_13_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_13_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_13_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_13_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_13_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_13_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_13_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_13_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_13_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_13_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_13_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_13_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_13_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_13_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_13_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_13_V_read[35]);
wire tmp_13_36;
assign tmp_13_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_13_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_13_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_13_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_13_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_13_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_13_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_13_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_13_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_13_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_13_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_13_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_13_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_13_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_13_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_13_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_13_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_13_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_13_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_13_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_13_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_13_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_13_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_13_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_13_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_13_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_13_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_13_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_13_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_13_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_13_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_13_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_13_V_read[36]);
wire tmp_13_37;
assign tmp_13_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_13_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_13_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_13_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_13_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_13_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_13_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_13_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_13_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_13_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_13_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_13_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_13_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_13_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_13_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_13_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_13_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_13_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_13_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_13_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_13_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_13_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_13_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_13_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_13_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_13_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_13_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_13_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_13_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_13_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_13_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_13_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_13_V_read[37]);
wire tmp_13_40;
assign tmp_13_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_13_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_13_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_13_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_13_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_13_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_13_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_13_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_13_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_13_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_13_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_13_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_13_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_13_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_13_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_13_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_13_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_13_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_13_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_13_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_13_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_13_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_13_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_13_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_13_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_13_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_13_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_13_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_13_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_13_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_13_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_13_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_13_V_read[40]);
wire tmp_13_41;
assign tmp_13_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_13_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_13_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_13_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_13_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_13_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_13_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_13_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_13_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_13_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_13_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_13_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_13_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_13_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_13_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_13_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_13_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_13_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_13_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_13_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_13_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_13_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_13_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_13_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_13_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_13_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_13_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_13_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_13_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_13_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_13_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_13_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_13_V_read[41]);
wire tmp_13_42;
assign tmp_13_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_13_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_13_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_13_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_13_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_13_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_13_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_13_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_13_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_13_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_13_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_13_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_13_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_13_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_13_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_13_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_13_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_13_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_13_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_13_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_13_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_13_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_13_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_13_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_13_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_13_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_13_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_13_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_13_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_13_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_13_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_13_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_13_V_read[42]);
wire tmp_13_43;
assign tmp_13_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_13_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_13_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_13_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_13_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_13_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_13_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_13_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_13_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_13_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_13_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_13_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_13_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_13_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_13_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_13_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_13_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_13_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_13_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_13_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_13_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_13_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_13_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_13_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_13_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_13_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_13_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_13_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_13_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_13_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_13_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_13_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_13_V_read[43]);
wire tmp_13_44;
assign tmp_13_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_13_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_13_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_13_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_13_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_13_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_13_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_13_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_13_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_13_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_13_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_13_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_13_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_13_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_13_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_13_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_13_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_13_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_13_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_13_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_13_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_13_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_13_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_13_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_13_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_13_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_13_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_13_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_13_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_13_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_13_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_13_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_13_V_read[44]);
wire tmp_13_45;
assign tmp_13_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_13_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_13_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_13_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_13_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_13_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_13_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_13_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_13_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_13_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_13_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_13_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_13_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_13_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_13_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_13_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_13_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_13_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_13_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_13_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_13_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_13_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_13_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_13_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_13_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_13_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_13_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_13_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_13_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_13_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_13_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_13_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_13_V_read[45]);
wire tmp_13_48;
assign tmp_13_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_13_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_13_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_13_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_13_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_13_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_13_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_13_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_13_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_13_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_13_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_13_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_13_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_13_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_13_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_13_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_13_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_13_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_13_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_13_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_13_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_13_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_13_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_13_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_13_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_13_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_13_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_13_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_13_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_13_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_13_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_13_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_13_V_read[48]);
wire tmp_13_49;
assign tmp_13_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_13_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_13_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_13_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_13_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_13_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_13_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_13_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_13_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_13_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_13_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_13_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_13_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_13_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_13_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_13_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_13_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_13_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_13_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_13_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_13_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_13_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_13_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_13_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_13_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_13_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_13_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_13_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_13_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_13_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_13_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_13_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_13_V_read[49]);
wire tmp_13_50;
assign tmp_13_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_13_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_13_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_13_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_13_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_13_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_13_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_13_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_13_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_13_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_13_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_13_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_13_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_13_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_13_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_13_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_13_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_13_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_13_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_13_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_13_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_13_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_13_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_13_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_13_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_13_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_13_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_13_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_13_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_13_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_13_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_13_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_13_V_read[50]);
wire tmp_13_51;
assign tmp_13_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_13_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_13_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_13_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_13_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_13_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_13_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_13_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_13_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_13_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_13_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_13_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_13_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_13_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_13_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_13_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_13_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_13_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_13_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_13_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_13_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_13_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_13_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_13_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_13_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_13_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_13_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_13_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_13_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_13_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_13_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_13_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_13_V_read[51]);
wire tmp_13_52;
assign tmp_13_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_13_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_13_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_13_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_13_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_13_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_13_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_13_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_13_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_13_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_13_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_13_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_13_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_13_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_13_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_13_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_13_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_13_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_13_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_13_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_13_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_13_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_13_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_13_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_13_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_13_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_13_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_13_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_13_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_13_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_13_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_13_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_13_V_read[52]);
wire tmp_13_53;
assign tmp_13_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_13_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_13_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_13_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_13_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_13_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_13_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_13_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_13_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_13_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_13_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_13_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_13_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_13_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_13_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_13_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_13_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_13_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_13_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_13_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_13_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_13_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_13_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_13_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_13_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_13_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_13_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_13_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_13_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_13_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_13_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_13_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_13_V_read[53]);
wire tmp_13_54;
assign tmp_13_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_13_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_13_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_13_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_13_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_13_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_13_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_13_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_13_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_13_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_13_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_13_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_13_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_13_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_13_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_13_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_13_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_13_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_13_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_13_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_13_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_13_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_13_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_13_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_13_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_13_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_13_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_13_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_13_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_13_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_13_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_13_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_13_V_read[54]);
wire tmp_13_55;
assign tmp_13_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_13_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_13_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_13_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_13_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_13_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_13_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_13_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_13_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_13_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_13_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_13_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_13_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_13_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_13_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_13_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_13_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_13_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_13_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_13_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_13_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_13_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_13_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_13_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_13_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_13_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_13_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_13_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_13_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_13_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_13_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_13_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_13_V_read[55]);
wire tmp_13_56;
assign tmp_13_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_13_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_13_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_13_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_13_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_13_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_13_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_13_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_13_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_13_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_13_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_13_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_13_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_13_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_13_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_13_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_13_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_13_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_13_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_13_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_13_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_13_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_13_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_13_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_13_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_13_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_13_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_13_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_13_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_13_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_13_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_13_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_13_V_read[56]);
wire tmp_13_57;
assign tmp_13_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_13_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_13_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_13_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_13_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_13_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_13_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_13_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_13_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_13_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_13_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_13_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_13_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_13_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_13_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_13_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_13_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_13_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_13_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_13_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_13_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_13_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_13_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_13_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_13_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_13_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_13_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_13_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_13_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_13_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_13_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_13_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_13_V_read[57]);
wire tmp_13_58;
assign tmp_13_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_13_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_13_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_13_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_13_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_13_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_13_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_13_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_13_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_13_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_13_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_13_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_13_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_13_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_13_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_13_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_13_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_13_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_13_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_13_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_13_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_13_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_13_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_13_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_13_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_13_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_13_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_13_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_13_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_13_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_13_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_13_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_13_V_read[58]);
wire tmp_13_59;
assign tmp_13_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_13_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_13_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_13_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_13_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_13_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_13_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_13_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_13_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_13_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_13_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_13_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_13_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_13_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_13_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_13_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_13_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_13_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_13_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_13_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_13_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_13_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_13_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_13_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_13_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_13_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_13_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_13_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_13_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_13_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_13_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_13_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_13_V_read[59]);
wire tmp_13_60;
assign tmp_13_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_13_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_13_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_13_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_13_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_13_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_13_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_13_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_13_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_13_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_13_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_13_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_13_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_13_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_13_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_13_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_13_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_13_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_13_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_13_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_13_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_13_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_13_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_13_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_13_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_13_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_13_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_13_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_13_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_13_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_13_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_13_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_13_V_read[60]);
wire tmp_13_61;
assign tmp_13_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_13_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_13_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_13_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_13_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_13_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_13_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_13_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_13_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_13_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_13_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_13_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_13_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_13_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_13_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_13_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_13_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_13_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_13_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_13_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_13_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_13_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_13_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_13_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_13_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_13_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_13_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_13_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_13_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_13_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_13_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_13_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_13_V_read[61]);
wire tmp_13_62;
assign tmp_13_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_13_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_13_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_13_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_13_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_13_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_13_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_13_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_13_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_13_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_13_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_13_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_13_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_13_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_13_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_13_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_13_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_13_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_13_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_13_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_13_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_13_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_13_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_13_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_13_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_13_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_13_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_13_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_13_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_13_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_13_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_13_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_13_V_read[62]);
wire tmp_13_63;
assign tmp_13_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_13_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_13_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_13_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_13_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_13_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_13_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_13_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_13_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_13_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_13_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_13_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_13_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_13_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_13_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_13_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_13_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_13_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_13_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_13_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_13_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_13_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_13_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_13_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_13_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_13_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_13_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_13_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_13_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_13_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_13_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_13_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_13_V_read[63]);
wire tmp_13_64;
assign tmp_13_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_13_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_13_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_13_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_13_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_13_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_13_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_13_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_13_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_13_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_13_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_13_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_13_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_13_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_13_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_13_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_13_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_13_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_13_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_13_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_13_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_13_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_13_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_13_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_13_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_13_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_13_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_13_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_13_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_13_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_13_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_13_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_13_V_read[64]);
wire tmp_13_65;
assign tmp_13_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_13_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_13_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_13_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_13_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_13_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_13_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_13_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_13_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_13_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_13_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_13_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_13_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_13_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_13_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_13_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_13_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_13_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_13_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_13_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_13_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_13_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_13_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_13_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_13_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_13_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_13_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_13_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_13_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_13_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_13_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_13_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_13_V_read[65]);
wire tmp_13_66;
assign tmp_13_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_13_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_13_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_13_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_13_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_13_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_13_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_13_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_13_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_13_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_13_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_13_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_13_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_13_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_13_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_13_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_13_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_13_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_13_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_13_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_13_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_13_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_13_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_13_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_13_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_13_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_13_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_13_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_13_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_13_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_13_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_13_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_13_V_read[66]);
wire tmp_13_67;
assign tmp_13_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_13_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_13_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_13_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_13_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_13_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_13_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_13_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_13_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_13_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_13_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_13_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_13_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_13_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_13_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_13_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_13_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_13_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_13_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_13_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_13_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_13_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_13_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_13_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_13_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_13_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_13_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_13_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_13_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_13_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_13_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_13_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_13_V_read[67]);
wire tmp_13_68;
assign tmp_13_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_13_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_13_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_13_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_13_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_13_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_13_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_13_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_13_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_13_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_13_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_13_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_13_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_13_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_13_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_13_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_13_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_13_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_13_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_13_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_13_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_13_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_13_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_13_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_13_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_13_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_13_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_13_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_13_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_13_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_13_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_13_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_13_V_read[68]);
wire tmp_13_70;
assign tmp_13_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_13_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_13_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_13_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_13_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_13_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_13_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_13_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_13_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_13_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_13_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_13_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_13_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_13_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_13_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_13_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_13_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_13_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_13_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_13_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_13_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_13_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_13_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_13_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_13_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_13_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_13_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_13_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_13_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_13_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_13_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_13_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_13_V_read[70]);
wire tmp_13_71;
assign tmp_13_71 = (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_13_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_13_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_13_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_13_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_13_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_13_V_read[71]) | (1 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_13_V_read[71]) | (0 &  in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_13_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_13_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_13_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_13_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_13_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_13_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_13_V_read[71]) | (1 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_13_V_read[71]) | (0 &  in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_13_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_13_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_13_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_13_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_13_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_13_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_13_V_read[71]) | (0 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_13_V_read[71]) | (1 & ~in_V[71] &  in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_13_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] &  weight_0_13_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] &  in_3_V[71] & ~weight_0_13_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] &  weight_0_13_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] &  in_2_V[71] & ~in_3_V[71] & ~weight_0_13_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] &  weight_0_13_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] &  in_3_V[71] & ~weight_0_13_V_read[71]) | (0 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] &  weight_0_13_V_read[71]) | (1 & ~in_V[71] & ~in_1_V[71] & ~in_2_V[71] & ~in_3_V[71] & ~weight_0_13_V_read[71]);
assign ap_return_13 = {tmp_13_0,tmp_13_1,tmp_13_2,tmp_13_3,tmp_13_4,tmp_13_5,1'b0,tmp_13_7,tmp_13_8,tmp_13_9,tmp_13_10,tmp_13_11,tmp_13_12,tmp_13_13,tmp_13_14,tmp_13_15,tmp_13_16,tmp_13_17,tmp_13_18,tmp_13_19,tmp_13_20,tmp_13_21,tmp_13_22,tmp_13_23,tmp_13_24,tmp_13_25,tmp_13_26,tmp_13_27,tmp_13_28,tmp_13_29,tmp_13_30,tmp_13_31,tmp_13_32,tmp_13_33,1'b0,tmp_13_35,tmp_13_36,tmp_13_37,1'b0,1'b0,tmp_13_40,tmp_13_41,tmp_13_42,tmp_13_43,tmp_13_44,tmp_13_45,1'b0,1'b0,tmp_13_48,tmp_13_49,tmp_13_50,tmp_13_51,tmp_13_52,tmp_13_53,tmp_13_54,tmp_13_55,tmp_13_56,tmp_13_57,tmp_13_58,tmp_13_59,tmp_13_60,tmp_13_61,tmp_13_62,tmp_13_63,tmp_13_64,tmp_13_65,tmp_13_66,tmp_13_67,tmp_13_68,1'b0,tmp_13_70,tmp_13_71};
wire tmp_14_0;
assign tmp_14_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_14_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_14_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_14_V_read[0]);
wire tmp_14_1;
assign tmp_14_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_14_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_14_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_14_V_read[1]);
wire tmp_14_2;
assign tmp_14_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_14_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_14_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_14_V_read[2]);
wire tmp_14_3;
assign tmp_14_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_14_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_14_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_14_V_read[3]);
wire tmp_14_4;
assign tmp_14_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_14_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_14_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_14_V_read[4]);
wire tmp_14_5;
assign tmp_14_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_14_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_14_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_14_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_14_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_14_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_14_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_14_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_14_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_14_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_14_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_14_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_14_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_14_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_14_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_14_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_14_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_14_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_14_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_14_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_14_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_14_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_14_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_14_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_14_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_14_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_14_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_14_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_14_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_14_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_14_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_14_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_14_V_read[5]);
wire tmp_14_6;
assign tmp_14_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_14_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_14_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_14_V_read[6]);
wire tmp_14_7;
assign tmp_14_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_14_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_14_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_14_V_read[7]);
wire tmp_14_8;
assign tmp_14_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_14_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_14_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_14_V_read[8]);
wire tmp_14_9;
assign tmp_14_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_14_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_14_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_14_V_read[9]);
wire tmp_14_10;
assign tmp_14_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_14_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_14_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_14_V_read[10]);
wire tmp_14_11;
assign tmp_14_11 = (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (1 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (1 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (0 &  in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] &  in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] &  in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] &  in_3_V[11] & ~weight_0_14_V_read[11]) | (0 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] &  weight_0_14_V_read[11]) | (1 & ~in_V[11] & ~in_1_V[11] & ~in_2_V[11] & ~in_3_V[11] & ~weight_0_14_V_read[11]);
wire tmp_14_12;
assign tmp_14_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_14_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_14_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_14_V_read[12]);
wire tmp_14_13;
assign tmp_14_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_14_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_14_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_14_V_read[13]);
wire tmp_14_15;
assign tmp_14_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_14_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_14_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_14_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_14_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_14_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_14_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_14_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_14_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_14_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_14_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_14_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_14_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_14_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_14_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_14_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_14_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_14_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_14_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_14_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_14_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_14_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_14_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_14_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_14_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_14_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_14_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_14_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_14_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_14_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_14_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_14_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_14_V_read[15]);
wire tmp_14_16;
assign tmp_14_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_14_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_14_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_14_V_read[16]);
wire tmp_14_17;
assign tmp_14_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_14_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_14_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_14_V_read[17]);
wire tmp_14_18;
assign tmp_14_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_14_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_14_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_14_V_read[18]);
wire tmp_14_19;
assign tmp_14_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_14_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_14_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_14_V_read[19]);
wire tmp_14_20;
assign tmp_14_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_14_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_14_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_14_V_read[20]);
wire tmp_14_21;
assign tmp_14_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_14_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_14_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_14_V_read[21]);
wire tmp_14_22;
assign tmp_14_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_14_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_14_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_14_V_read[22]);
wire tmp_14_23;
assign tmp_14_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_14_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_14_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_14_V_read[23]);
wire tmp_14_24;
assign tmp_14_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_14_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_14_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_14_V_read[24]);
wire tmp_14_25;
assign tmp_14_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_14_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_14_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_14_V_read[25]);
wire tmp_14_26;
assign tmp_14_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_14_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_14_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_14_V_read[26]);
wire tmp_14_27;
assign tmp_14_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_14_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_14_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_14_V_read[27]);
wire tmp_14_28;
assign tmp_14_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_14_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_14_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_14_V_read[28]);
wire tmp_14_29;
assign tmp_14_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_14_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_14_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_14_V_read[29]);
wire tmp_14_30;
assign tmp_14_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_14_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_14_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_14_V_read[30]);
wire tmp_14_32;
assign tmp_14_32 = (1 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_14_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_14_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_14_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_14_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_14_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_14_V_read[32]) | (1 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_14_V_read[32]) | (0 &  in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_14_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_14_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_14_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_14_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_14_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_14_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_14_V_read[32]) | (1 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_14_V_read[32]) | (0 &  in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_14_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_14_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_14_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_14_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_14_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_14_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_14_V_read[32]) | (0 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_14_V_read[32]) | (1 & ~in_V[32] &  in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_14_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] &  weight_0_14_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] &  in_3_V[32] & ~weight_0_14_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] &  weight_0_14_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] &  in_2_V[32] & ~in_3_V[32] & ~weight_0_14_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] &  weight_0_14_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] &  in_3_V[32] & ~weight_0_14_V_read[32]) | (0 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] &  weight_0_14_V_read[32]) | (1 & ~in_V[32] & ~in_1_V[32] & ~in_2_V[32] & ~in_3_V[32] & ~weight_0_14_V_read[32]);
wire tmp_14_33;
assign tmp_14_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_14_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_14_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_14_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_14_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_14_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_14_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_14_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_14_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_14_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_14_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_14_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_14_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_14_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_14_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_14_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_14_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_14_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_14_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_14_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_14_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_14_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_14_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_14_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_14_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_14_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_14_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_14_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_14_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_14_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_14_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_14_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_14_V_read[33]);
wire tmp_14_34;
assign tmp_14_34 = (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_14_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_14_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_14_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_14_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_14_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_14_V_read[34]) | (1 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_14_V_read[34]) | (0 &  in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_14_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_14_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_14_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_14_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_14_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_14_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_14_V_read[34]) | (1 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_14_V_read[34]) | (0 &  in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_14_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_14_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_14_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_14_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_14_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_14_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_14_V_read[34]) | (0 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_14_V_read[34]) | (1 & ~in_V[34] &  in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_14_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] &  weight_0_14_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] &  in_3_V[34] & ~weight_0_14_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] &  weight_0_14_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] &  in_2_V[34] & ~in_3_V[34] & ~weight_0_14_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] &  weight_0_14_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] &  in_3_V[34] & ~weight_0_14_V_read[34]) | (0 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] &  weight_0_14_V_read[34]) | (1 & ~in_V[34] & ~in_1_V[34] & ~in_2_V[34] & ~in_3_V[34] & ~weight_0_14_V_read[34]);
wire tmp_14_35;
assign tmp_14_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_14_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_14_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_14_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_14_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_14_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_14_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_14_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_14_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_14_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_14_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_14_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_14_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_14_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_14_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_14_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_14_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_14_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_14_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_14_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_14_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_14_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_14_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_14_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_14_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_14_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_14_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_14_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_14_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_14_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_14_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_14_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_14_V_read[35]);
wire tmp_14_36;
assign tmp_14_36 = (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_14_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_14_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_14_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_14_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_14_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_14_V_read[36]) | (1 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_14_V_read[36]) | (0 &  in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_14_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_14_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_14_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_14_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_14_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_14_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_14_V_read[36]) | (1 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_14_V_read[36]) | (0 &  in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_14_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_14_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_14_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_14_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_14_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_14_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_14_V_read[36]) | (0 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_14_V_read[36]) | (1 & ~in_V[36] &  in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_14_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] &  weight_0_14_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] &  in_3_V[36] & ~weight_0_14_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] &  weight_0_14_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] &  in_2_V[36] & ~in_3_V[36] & ~weight_0_14_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] &  weight_0_14_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] &  in_3_V[36] & ~weight_0_14_V_read[36]) | (0 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] &  weight_0_14_V_read[36]) | (1 & ~in_V[36] & ~in_1_V[36] & ~in_2_V[36] & ~in_3_V[36] & ~weight_0_14_V_read[36]);
wire tmp_14_38;
assign tmp_14_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_14_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_14_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_14_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_14_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_14_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_14_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_14_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_14_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_14_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_14_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_14_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_14_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_14_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_14_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_14_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_14_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_14_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_14_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_14_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_14_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_14_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_14_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_14_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_14_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_14_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_14_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_14_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_14_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_14_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_14_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_14_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_14_V_read[38]);
wire tmp_14_39;
assign tmp_14_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_14_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_14_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_14_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_14_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_14_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_14_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_14_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_14_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_14_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_14_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_14_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_14_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_14_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_14_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_14_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_14_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_14_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_14_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_14_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_14_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_14_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_14_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_14_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_14_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_14_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_14_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_14_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_14_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_14_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_14_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_14_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_14_V_read[39]);
wire tmp_14_40;
assign tmp_14_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_14_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_14_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_14_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_14_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_14_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_14_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_14_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_14_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_14_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_14_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_14_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_14_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_14_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_14_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_14_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_14_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_14_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_14_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_14_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_14_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_14_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_14_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_14_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_14_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_14_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_14_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_14_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_14_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_14_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_14_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_14_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_14_V_read[40]);
wire tmp_14_41;
assign tmp_14_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_14_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_14_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_14_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_14_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_14_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_14_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_14_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_14_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_14_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_14_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_14_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_14_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_14_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_14_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_14_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_14_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_14_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_14_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_14_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_14_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_14_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_14_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_14_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_14_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_14_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_14_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_14_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_14_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_14_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_14_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_14_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_14_V_read[41]);
wire tmp_14_42;
assign tmp_14_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_14_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_14_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_14_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_14_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_14_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_14_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_14_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_14_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_14_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_14_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_14_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_14_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_14_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_14_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_14_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_14_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_14_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_14_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_14_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_14_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_14_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_14_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_14_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_14_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_14_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_14_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_14_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_14_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_14_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_14_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_14_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_14_V_read[42]);
wire tmp_14_43;
assign tmp_14_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_14_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_14_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_14_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_14_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_14_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_14_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_14_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_14_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_14_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_14_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_14_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_14_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_14_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_14_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_14_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_14_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_14_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_14_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_14_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_14_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_14_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_14_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_14_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_14_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_14_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_14_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_14_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_14_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_14_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_14_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_14_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_14_V_read[43]);
wire tmp_14_44;
assign tmp_14_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_14_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_14_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_14_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_14_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_14_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_14_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_14_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_14_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_14_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_14_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_14_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_14_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_14_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_14_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_14_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_14_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_14_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_14_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_14_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_14_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_14_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_14_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_14_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_14_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_14_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_14_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_14_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_14_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_14_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_14_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_14_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_14_V_read[44]);
wire tmp_14_45;
assign tmp_14_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_14_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_14_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_14_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_14_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_14_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_14_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_14_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_14_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_14_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_14_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_14_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_14_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_14_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_14_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_14_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_14_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_14_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_14_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_14_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_14_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_14_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_14_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_14_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_14_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_14_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_14_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_14_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_14_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_14_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_14_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_14_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_14_V_read[45]);
wire tmp_14_46;
assign tmp_14_46 = (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_14_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_14_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_14_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_14_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_14_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_14_V_read[46]) | (1 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_14_V_read[46]) | (0 &  in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_14_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_14_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_14_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_14_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_14_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_14_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_14_V_read[46]) | (1 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_14_V_read[46]) | (0 &  in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_14_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_14_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_14_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_14_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_14_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_14_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_14_V_read[46]) | (0 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_14_V_read[46]) | (1 & ~in_V[46] &  in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_14_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] &  weight_0_14_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] &  in_3_V[46] & ~weight_0_14_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] &  weight_0_14_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] &  in_2_V[46] & ~in_3_V[46] & ~weight_0_14_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] &  weight_0_14_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] &  in_3_V[46] & ~weight_0_14_V_read[46]) | (0 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] &  weight_0_14_V_read[46]) | (1 & ~in_V[46] & ~in_1_V[46] & ~in_2_V[46] & ~in_3_V[46] & ~weight_0_14_V_read[46]);
wire tmp_14_47;
assign tmp_14_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_14_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_14_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_14_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_14_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_14_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_14_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_14_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_14_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_14_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_14_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_14_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_14_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_14_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_14_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_14_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_14_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_14_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_14_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_14_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_14_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_14_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_14_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_14_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_14_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_14_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_14_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_14_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_14_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_14_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_14_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_14_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_14_V_read[47]);
wire tmp_14_48;
assign tmp_14_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_14_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_14_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_14_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_14_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_14_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_14_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_14_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_14_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_14_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_14_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_14_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_14_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_14_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_14_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_14_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_14_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_14_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_14_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_14_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_14_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_14_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_14_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_14_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_14_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_14_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_14_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_14_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_14_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_14_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_14_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_14_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_14_V_read[48]);
wire tmp_14_49;
assign tmp_14_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_14_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_14_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_14_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_14_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_14_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_14_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_14_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_14_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_14_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_14_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_14_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_14_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_14_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_14_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_14_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_14_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_14_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_14_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_14_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_14_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_14_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_14_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_14_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_14_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_14_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_14_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_14_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_14_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_14_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_14_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_14_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_14_V_read[49]);
wire tmp_14_50;
assign tmp_14_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_14_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_14_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_14_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_14_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_14_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_14_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_14_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_14_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_14_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_14_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_14_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_14_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_14_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_14_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_14_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_14_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_14_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_14_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_14_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_14_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_14_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_14_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_14_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_14_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_14_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_14_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_14_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_14_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_14_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_14_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_14_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_14_V_read[50]);
wire tmp_14_51;
assign tmp_14_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_14_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_14_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_14_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_14_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_14_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_14_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_14_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_14_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_14_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_14_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_14_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_14_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_14_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_14_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_14_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_14_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_14_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_14_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_14_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_14_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_14_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_14_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_14_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_14_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_14_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_14_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_14_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_14_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_14_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_14_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_14_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_14_V_read[51]);
wire tmp_14_52;
assign tmp_14_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_14_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_14_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_14_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_14_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_14_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_14_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_14_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_14_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_14_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_14_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_14_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_14_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_14_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_14_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_14_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_14_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_14_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_14_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_14_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_14_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_14_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_14_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_14_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_14_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_14_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_14_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_14_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_14_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_14_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_14_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_14_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_14_V_read[52]);
wire tmp_14_53;
assign tmp_14_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_14_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_14_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_14_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_14_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_14_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_14_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_14_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_14_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_14_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_14_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_14_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_14_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_14_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_14_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_14_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_14_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_14_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_14_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_14_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_14_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_14_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_14_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_14_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_14_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_14_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_14_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_14_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_14_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_14_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_14_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_14_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_14_V_read[53]);
wire tmp_14_54;
assign tmp_14_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_14_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_14_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_14_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_14_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_14_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_14_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_14_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_14_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_14_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_14_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_14_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_14_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_14_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_14_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_14_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_14_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_14_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_14_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_14_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_14_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_14_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_14_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_14_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_14_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_14_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_14_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_14_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_14_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_14_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_14_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_14_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_14_V_read[54]);
wire tmp_14_55;
assign tmp_14_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_14_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_14_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_14_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_14_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_14_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_14_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_14_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_14_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_14_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_14_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_14_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_14_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_14_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_14_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_14_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_14_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_14_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_14_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_14_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_14_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_14_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_14_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_14_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_14_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_14_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_14_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_14_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_14_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_14_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_14_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_14_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_14_V_read[55]);
wire tmp_14_56;
assign tmp_14_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_14_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_14_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_14_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_14_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_14_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_14_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_14_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_14_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_14_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_14_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_14_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_14_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_14_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_14_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_14_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_14_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_14_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_14_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_14_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_14_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_14_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_14_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_14_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_14_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_14_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_14_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_14_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_14_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_14_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_14_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_14_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_14_V_read[56]);
wire tmp_14_57;
assign tmp_14_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_14_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_14_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_14_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_14_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_14_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_14_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_14_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_14_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_14_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_14_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_14_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_14_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_14_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_14_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_14_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_14_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_14_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_14_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_14_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_14_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_14_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_14_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_14_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_14_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_14_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_14_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_14_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_14_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_14_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_14_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_14_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_14_V_read[57]);
wire tmp_14_58;
assign tmp_14_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_14_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_14_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_14_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_14_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_14_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_14_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_14_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_14_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_14_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_14_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_14_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_14_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_14_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_14_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_14_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_14_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_14_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_14_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_14_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_14_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_14_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_14_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_14_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_14_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_14_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_14_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_14_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_14_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_14_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_14_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_14_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_14_V_read[58]);
wire tmp_14_59;
assign tmp_14_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_14_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_14_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_14_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_14_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_14_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_14_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_14_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_14_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_14_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_14_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_14_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_14_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_14_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_14_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_14_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_14_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_14_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_14_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_14_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_14_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_14_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_14_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_14_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_14_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_14_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_14_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_14_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_14_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_14_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_14_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_14_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_14_V_read[59]);
wire tmp_14_61;
assign tmp_14_61 = (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_14_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_14_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_14_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_14_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_14_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_14_V_read[61]) | (1 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_14_V_read[61]) | (0 &  in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_14_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_14_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_14_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_14_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_14_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_14_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_14_V_read[61]) | (1 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_14_V_read[61]) | (0 &  in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_14_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_14_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_14_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_14_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_14_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_14_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_14_V_read[61]) | (0 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_14_V_read[61]) | (1 & ~in_V[61] &  in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_14_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] &  weight_0_14_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] &  in_3_V[61] & ~weight_0_14_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] &  weight_0_14_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] &  in_2_V[61] & ~in_3_V[61] & ~weight_0_14_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] &  weight_0_14_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] &  in_3_V[61] & ~weight_0_14_V_read[61]) | (0 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] &  weight_0_14_V_read[61]) | (1 & ~in_V[61] & ~in_1_V[61] & ~in_2_V[61] & ~in_3_V[61] & ~weight_0_14_V_read[61]);
wire tmp_14_64;
assign tmp_14_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_14_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_14_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_14_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_14_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_14_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_14_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_14_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_14_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_14_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_14_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_14_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_14_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_14_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_14_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_14_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_14_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_14_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_14_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_14_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_14_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_14_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_14_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_14_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_14_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_14_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_14_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_14_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_14_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_14_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_14_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_14_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_14_V_read[64]);
wire tmp_14_65;
assign tmp_14_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_14_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_14_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_14_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_14_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_14_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_14_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_14_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_14_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_14_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_14_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_14_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_14_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_14_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_14_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_14_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_14_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_14_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_14_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_14_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_14_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_14_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_14_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_14_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_14_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_14_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_14_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_14_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_14_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_14_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_14_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_14_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_14_V_read[65]);
wire tmp_14_66;
assign tmp_14_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_14_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_14_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_14_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_14_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_14_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_14_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_14_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_14_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_14_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_14_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_14_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_14_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_14_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_14_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_14_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_14_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_14_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_14_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_14_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_14_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_14_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_14_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_14_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_14_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_14_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_14_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_14_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_14_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_14_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_14_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_14_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_14_V_read[66]);
wire tmp_14_67;
assign tmp_14_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_14_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_14_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_14_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_14_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_14_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_14_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_14_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_14_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_14_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_14_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_14_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_14_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_14_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_14_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_14_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_14_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_14_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_14_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_14_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_14_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_14_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_14_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_14_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_14_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_14_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_14_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_14_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_14_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_14_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_14_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_14_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_14_V_read[67]);
wire tmp_14_69;
assign tmp_14_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_14_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_14_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_14_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_14_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_14_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_14_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_14_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_14_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_14_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_14_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_14_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_14_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_14_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_14_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_14_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_14_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_14_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_14_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_14_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_14_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_14_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_14_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_14_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_14_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_14_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_14_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_14_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_14_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_14_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_14_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_14_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_14_V_read[69]);
wire tmp_14_70;
assign tmp_14_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_14_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_14_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_14_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_14_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_14_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_14_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_14_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_14_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_14_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_14_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_14_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_14_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_14_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_14_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_14_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_14_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_14_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_14_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_14_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_14_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_14_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_14_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_14_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_14_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_14_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_14_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_14_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_14_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_14_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_14_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_14_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_14_V_read[70]);
assign ap_return_14 = {tmp_14_0,tmp_14_1,tmp_14_2,tmp_14_3,tmp_14_4,tmp_14_5,tmp_14_6,tmp_14_7,tmp_14_8,tmp_14_9,tmp_14_10,tmp_14_11,tmp_14_12,tmp_14_13,1'b0,tmp_14_15,tmp_14_16,tmp_14_17,tmp_14_18,tmp_14_19,tmp_14_20,tmp_14_21,tmp_14_22,tmp_14_23,tmp_14_24,tmp_14_25,tmp_14_26,tmp_14_27,tmp_14_28,tmp_14_29,tmp_14_30,1'b0,tmp_14_32,tmp_14_33,tmp_14_34,tmp_14_35,tmp_14_36,1'b0,tmp_14_38,tmp_14_39,tmp_14_40,tmp_14_41,tmp_14_42,tmp_14_43,tmp_14_44,tmp_14_45,tmp_14_46,tmp_14_47,tmp_14_48,tmp_14_49,tmp_14_50,tmp_14_51,tmp_14_52,tmp_14_53,tmp_14_54,tmp_14_55,tmp_14_56,tmp_14_57,tmp_14_58,tmp_14_59,1'b0,tmp_14_61,1'b0,1'b0,tmp_14_64,tmp_14_65,tmp_14_66,tmp_14_67,1'b0,tmp_14_69,tmp_14_70,1'b0};
wire tmp_15_0;
assign tmp_15_0 = (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (1 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (1 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (0 &  in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] &  in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] &  in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] &  in_3_V[0] & ~weight_0_15_V_read[0]) | (0 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] &  weight_0_15_V_read[0]) | (1 & ~in_V[0] & ~in_1_V[0] & ~in_2_V[0] & ~in_3_V[0] & ~weight_0_15_V_read[0]);
wire tmp_15_1;
assign tmp_15_1 = (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (1 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (1 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (0 &  in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] &  in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] &  in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] &  in_3_V[1] & ~weight_0_15_V_read[1]) | (0 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] &  weight_0_15_V_read[1]) | (1 & ~in_V[1] & ~in_1_V[1] & ~in_2_V[1] & ~in_3_V[1] & ~weight_0_15_V_read[1]);
wire tmp_15_2;
assign tmp_15_2 = (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (1 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (1 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (0 &  in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] &  in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] &  in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] &  in_3_V[2] & ~weight_0_15_V_read[2]) | (0 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] &  weight_0_15_V_read[2]) | (1 & ~in_V[2] & ~in_1_V[2] & ~in_2_V[2] & ~in_3_V[2] & ~weight_0_15_V_read[2]);
wire tmp_15_3;
assign tmp_15_3 = (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (1 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (0 &  in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] &  in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] &  in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] &  in_3_V[3] & ~weight_0_15_V_read[3]) | (0 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] &  weight_0_15_V_read[3]) | (1 & ~in_V[3] & ~in_1_V[3] & ~in_2_V[3] & ~in_3_V[3] & ~weight_0_15_V_read[3]);
wire tmp_15_4;
assign tmp_15_4 = (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (1 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (1 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (0 &  in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] &  in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] &  in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] &  in_3_V[4] & ~weight_0_15_V_read[4]) | (0 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] &  weight_0_15_V_read[4]) | (1 & ~in_V[4] & ~in_1_V[4] & ~in_2_V[4] & ~in_3_V[4] & ~weight_0_15_V_read[4]);
wire tmp_15_5;
assign tmp_15_5 = (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (1 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (1 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (0 &  in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] &  in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] &  in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] &  in_3_V[5] & ~weight_0_15_V_read[5]) | (0 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] &  weight_0_15_V_read[5]) | (1 & ~in_V[5] & ~in_1_V[5] & ~in_2_V[5] & ~in_3_V[5] & ~weight_0_15_V_read[5]);
wire tmp_15_6;
assign tmp_15_6 = (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (1 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (1 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (0 &  in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] &  in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] &  in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] &  in_3_V[6] & ~weight_0_15_V_read[6]) | (0 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] &  weight_0_15_V_read[6]) | (1 & ~in_V[6] & ~in_1_V[6] & ~in_2_V[6] & ~in_3_V[6] & ~weight_0_15_V_read[6]);
wire tmp_15_7;
assign tmp_15_7 = (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (1 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (0 &  in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] &  in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] &  in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] &  in_3_V[7] & ~weight_0_15_V_read[7]) | (0 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] &  weight_0_15_V_read[7]) | (1 & ~in_V[7] & ~in_1_V[7] & ~in_2_V[7] & ~in_3_V[7] & ~weight_0_15_V_read[7]);
wire tmp_15_8;
assign tmp_15_8 = (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (1 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (1 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (0 &  in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] &  in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] &  in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] &  in_3_V[8] & ~weight_0_15_V_read[8]) | (0 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] &  weight_0_15_V_read[8]) | (1 & ~in_V[8] & ~in_1_V[8] & ~in_2_V[8] & ~in_3_V[8] & ~weight_0_15_V_read[8]);
wire tmp_15_9;
assign tmp_15_9 = (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (1 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (0 &  in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] &  in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] &  in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] &  in_3_V[9] & ~weight_0_15_V_read[9]) | (0 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] &  weight_0_15_V_read[9]) | (1 & ~in_V[9] & ~in_1_V[9] & ~in_2_V[9] & ~in_3_V[9] & ~weight_0_15_V_read[9]);
wire tmp_15_10;
assign tmp_15_10 = (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (1 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (1 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (0 &  in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] &  in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] &  in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] &  in_3_V[10] & ~weight_0_15_V_read[10]) | (0 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] &  weight_0_15_V_read[10]) | (1 & ~in_V[10] & ~in_1_V[10] & ~in_2_V[10] & ~in_3_V[10] & ~weight_0_15_V_read[10]);
wire tmp_15_12;
assign tmp_15_12 = (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (1 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (1 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (0 &  in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] &  in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] &  in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] &  in_3_V[12] & ~weight_0_15_V_read[12]) | (0 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] &  weight_0_15_V_read[12]) | (1 & ~in_V[12] & ~in_1_V[12] & ~in_2_V[12] & ~in_3_V[12] & ~weight_0_15_V_read[12]);
wire tmp_15_13;
assign tmp_15_13 = (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (1 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (1 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (0 &  in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] &  in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] &  in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] &  in_3_V[13] & ~weight_0_15_V_read[13]) | (0 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] &  weight_0_15_V_read[13]) | (1 & ~in_V[13] & ~in_1_V[13] & ~in_2_V[13] & ~in_3_V[13] & ~weight_0_15_V_read[13]);
wire tmp_15_14;
assign tmp_15_14 = (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (1 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (1 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (0 &  in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] &  in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] &  in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] &  in_3_V[14] & ~weight_0_15_V_read[14]) | (0 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] &  weight_0_15_V_read[14]) | (1 & ~in_V[14] & ~in_1_V[14] & ~in_2_V[14] & ~in_3_V[14] & ~weight_0_15_V_read[14]);
wire tmp_15_15;
assign tmp_15_15 = (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (1 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (1 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (0 &  in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] &  in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] &  in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] &  in_3_V[15] & ~weight_0_15_V_read[15]) | (0 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] &  weight_0_15_V_read[15]) | (1 & ~in_V[15] & ~in_1_V[15] & ~in_2_V[15] & ~in_3_V[15] & ~weight_0_15_V_read[15]);
wire tmp_15_16;
assign tmp_15_16 = (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (1 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (1 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (0 &  in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] &  in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] &  in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] &  in_3_V[16] & ~weight_0_15_V_read[16]) | (0 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] &  weight_0_15_V_read[16]) | (1 & ~in_V[16] & ~in_1_V[16] & ~in_2_V[16] & ~in_3_V[16] & ~weight_0_15_V_read[16]);
wire tmp_15_17;
assign tmp_15_17 = (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (1 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (1 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (0 &  in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] &  in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] &  in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] &  in_3_V[17] & ~weight_0_15_V_read[17]) | (0 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] &  weight_0_15_V_read[17]) | (1 & ~in_V[17] & ~in_1_V[17] & ~in_2_V[17] & ~in_3_V[17] & ~weight_0_15_V_read[17]);
wire tmp_15_18;
assign tmp_15_18 = (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (1 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (0 &  in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] &  in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] &  in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] &  in_3_V[18] & ~weight_0_15_V_read[18]) | (0 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] &  weight_0_15_V_read[18]) | (1 & ~in_V[18] & ~in_1_V[18] & ~in_2_V[18] & ~in_3_V[18] & ~weight_0_15_V_read[18]);
wire tmp_15_19;
assign tmp_15_19 = (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (1 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (0 &  in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] &  in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] &  in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] &  in_3_V[19] & ~weight_0_15_V_read[19]) | (0 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] &  weight_0_15_V_read[19]) | (1 & ~in_V[19] & ~in_1_V[19] & ~in_2_V[19] & ~in_3_V[19] & ~weight_0_15_V_read[19]);
wire tmp_15_20;
assign tmp_15_20 = (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (1 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (0 &  in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] &  in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] &  in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] &  in_3_V[20] & ~weight_0_15_V_read[20]) | (0 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] &  weight_0_15_V_read[20]) | (1 & ~in_V[20] & ~in_1_V[20] & ~in_2_V[20] & ~in_3_V[20] & ~weight_0_15_V_read[20]);
wire tmp_15_21;
assign tmp_15_21 = (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (1 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (0 &  in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] &  in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] &  in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] &  in_3_V[21] & ~weight_0_15_V_read[21]) | (0 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] &  weight_0_15_V_read[21]) | (1 & ~in_V[21] & ~in_1_V[21] & ~in_2_V[21] & ~in_3_V[21] & ~weight_0_15_V_read[21]);
wire tmp_15_22;
assign tmp_15_22 = (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (1 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (1 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (0 &  in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] &  in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] &  in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] &  in_3_V[22] & ~weight_0_15_V_read[22]) | (0 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] &  weight_0_15_V_read[22]) | (1 & ~in_V[22] & ~in_1_V[22] & ~in_2_V[22] & ~in_3_V[22] & ~weight_0_15_V_read[22]);
wire tmp_15_23;
assign tmp_15_23 = (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (1 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (0 &  in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] &  in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] &  in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] &  in_3_V[23] & ~weight_0_15_V_read[23]) | (0 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] &  weight_0_15_V_read[23]) | (1 & ~in_V[23] & ~in_1_V[23] & ~in_2_V[23] & ~in_3_V[23] & ~weight_0_15_V_read[23]);
wire tmp_15_24;
assign tmp_15_24 = (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (1 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (1 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (0 &  in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] &  in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] &  in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] &  in_3_V[24] & ~weight_0_15_V_read[24]) | (0 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] &  weight_0_15_V_read[24]) | (1 & ~in_V[24] & ~in_1_V[24] & ~in_2_V[24] & ~in_3_V[24] & ~weight_0_15_V_read[24]);
wire tmp_15_25;
assign tmp_15_25 = (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (1 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (1 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (0 &  in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] &  in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] &  in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] &  in_3_V[25] & ~weight_0_15_V_read[25]) | (0 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] &  weight_0_15_V_read[25]) | (1 & ~in_V[25] & ~in_1_V[25] & ~in_2_V[25] & ~in_3_V[25] & ~weight_0_15_V_read[25]);
wire tmp_15_26;
assign tmp_15_26 = (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (1 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (1 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (0 &  in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] &  in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] &  in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] &  in_3_V[26] & ~weight_0_15_V_read[26]) | (0 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] &  weight_0_15_V_read[26]) | (1 & ~in_V[26] & ~in_1_V[26] & ~in_2_V[26] & ~in_3_V[26] & ~weight_0_15_V_read[26]);
wire tmp_15_27;
assign tmp_15_27 = (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (1 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (1 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (0 &  in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] &  in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] &  in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] &  in_3_V[27] & ~weight_0_15_V_read[27]) | (0 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] &  weight_0_15_V_read[27]) | (1 & ~in_V[27] & ~in_1_V[27] & ~in_2_V[27] & ~in_3_V[27] & ~weight_0_15_V_read[27]);
wire tmp_15_28;
assign tmp_15_28 = (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (1 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (1 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (0 &  in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] &  in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] &  in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] &  in_3_V[28] & ~weight_0_15_V_read[28]) | (0 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] &  weight_0_15_V_read[28]) | (1 & ~in_V[28] & ~in_1_V[28] & ~in_2_V[28] & ~in_3_V[28] & ~weight_0_15_V_read[28]);
wire tmp_15_29;
assign tmp_15_29 = (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (1 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (0 &  in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] &  in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] &  in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] &  in_3_V[29] & ~weight_0_15_V_read[29]) | (0 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] &  weight_0_15_V_read[29]) | (1 & ~in_V[29] & ~in_1_V[29] & ~in_2_V[29] & ~in_3_V[29] & ~weight_0_15_V_read[29]);
wire tmp_15_30;
assign tmp_15_30 = (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (1 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (1 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (0 &  in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] &  in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] &  in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] &  in_3_V[30] & ~weight_0_15_V_read[30]) | (0 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] &  weight_0_15_V_read[30]) | (1 & ~in_V[30] & ~in_1_V[30] & ~in_2_V[30] & ~in_3_V[30] & ~weight_0_15_V_read[30]);
wire tmp_15_33;
assign tmp_15_33 = (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_15_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_15_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_15_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_15_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_15_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_15_V_read[33]) | (1 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_15_V_read[33]) | (0 &  in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_15_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_15_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_15_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_15_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_15_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_15_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_15_V_read[33]) | (1 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_15_V_read[33]) | (0 &  in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_15_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_15_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_15_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_15_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_15_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_15_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_15_V_read[33]) | (0 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_15_V_read[33]) | (1 & ~in_V[33] &  in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_15_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] &  weight_0_15_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] &  in_3_V[33] & ~weight_0_15_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] &  weight_0_15_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] &  in_2_V[33] & ~in_3_V[33] & ~weight_0_15_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] &  weight_0_15_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] &  in_3_V[33] & ~weight_0_15_V_read[33]) | (0 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] &  weight_0_15_V_read[33]) | (1 & ~in_V[33] & ~in_1_V[33] & ~in_2_V[33] & ~in_3_V[33] & ~weight_0_15_V_read[33]);
wire tmp_15_35;
assign tmp_15_35 = (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_15_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_15_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_15_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_15_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_15_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_15_V_read[35]) | (1 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_15_V_read[35]) | (0 &  in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_15_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_15_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_15_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_15_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_15_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_15_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_15_V_read[35]) | (1 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_15_V_read[35]) | (0 &  in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_15_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_15_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_15_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_15_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_15_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_15_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_15_V_read[35]) | (0 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_15_V_read[35]) | (1 & ~in_V[35] &  in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_15_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] &  weight_0_15_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] &  in_3_V[35] & ~weight_0_15_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] &  weight_0_15_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] &  in_2_V[35] & ~in_3_V[35] & ~weight_0_15_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] &  weight_0_15_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] &  in_3_V[35] & ~weight_0_15_V_read[35]) | (0 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] &  weight_0_15_V_read[35]) | (1 & ~in_V[35] & ~in_1_V[35] & ~in_2_V[35] & ~in_3_V[35] & ~weight_0_15_V_read[35]);
wire tmp_15_37;
assign tmp_15_37 = (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_15_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_15_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_15_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_15_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_15_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_15_V_read[37]) | (1 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_15_V_read[37]) | (0 &  in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_15_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_15_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_15_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_15_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_15_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_15_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_15_V_read[37]) | (1 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_15_V_read[37]) | (0 &  in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_15_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_15_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_15_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_15_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_15_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_15_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_15_V_read[37]) | (0 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_15_V_read[37]) | (1 & ~in_V[37] &  in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_15_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] &  weight_0_15_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] &  in_3_V[37] & ~weight_0_15_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] &  weight_0_15_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] &  in_2_V[37] & ~in_3_V[37] & ~weight_0_15_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] &  weight_0_15_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] &  in_3_V[37] & ~weight_0_15_V_read[37]) | (0 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] &  weight_0_15_V_read[37]) | (1 & ~in_V[37] & ~in_1_V[37] & ~in_2_V[37] & ~in_3_V[37] & ~weight_0_15_V_read[37]);
wire tmp_15_38;
assign tmp_15_38 = (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_15_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_15_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_15_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_15_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_15_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_15_V_read[38]) | (1 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_15_V_read[38]) | (0 &  in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_15_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_15_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_15_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_15_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_15_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_15_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_15_V_read[38]) | (1 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_15_V_read[38]) | (0 &  in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_15_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_15_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_15_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_15_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_15_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_15_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_15_V_read[38]) | (0 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_15_V_read[38]) | (1 & ~in_V[38] &  in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_15_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] &  weight_0_15_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] &  in_3_V[38] & ~weight_0_15_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] &  weight_0_15_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] &  in_2_V[38] & ~in_3_V[38] & ~weight_0_15_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] &  weight_0_15_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] &  in_3_V[38] & ~weight_0_15_V_read[38]) | (0 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] &  weight_0_15_V_read[38]) | (1 & ~in_V[38] & ~in_1_V[38] & ~in_2_V[38] & ~in_3_V[38] & ~weight_0_15_V_read[38]);
wire tmp_15_39;
assign tmp_15_39 = (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_15_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_15_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_15_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_15_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_15_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_15_V_read[39]) | (1 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_15_V_read[39]) | (0 &  in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_15_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_15_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_15_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_15_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_15_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_15_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_15_V_read[39]) | (1 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_15_V_read[39]) | (0 &  in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_15_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_15_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_15_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_15_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_15_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_15_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_15_V_read[39]) | (0 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_15_V_read[39]) | (1 & ~in_V[39] &  in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_15_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] &  weight_0_15_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] &  in_3_V[39] & ~weight_0_15_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] &  weight_0_15_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] &  in_2_V[39] & ~in_3_V[39] & ~weight_0_15_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] &  weight_0_15_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] &  in_3_V[39] & ~weight_0_15_V_read[39]) | (0 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] &  weight_0_15_V_read[39]) | (1 & ~in_V[39] & ~in_1_V[39] & ~in_2_V[39] & ~in_3_V[39] & ~weight_0_15_V_read[39]);
wire tmp_15_40;
assign tmp_15_40 = (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_15_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_15_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_15_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_15_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_15_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_15_V_read[40]) | (1 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_15_V_read[40]) | (0 &  in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_15_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_15_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_15_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_15_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_15_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_15_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_15_V_read[40]) | (1 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_15_V_read[40]) | (0 &  in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_15_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_15_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_15_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_15_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_15_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_15_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_15_V_read[40]) | (0 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_15_V_read[40]) | (1 & ~in_V[40] &  in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_15_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] &  weight_0_15_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] &  in_3_V[40] & ~weight_0_15_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] &  weight_0_15_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] &  in_2_V[40] & ~in_3_V[40] & ~weight_0_15_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] &  weight_0_15_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] &  in_3_V[40] & ~weight_0_15_V_read[40]) | (0 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] &  weight_0_15_V_read[40]) | (1 & ~in_V[40] & ~in_1_V[40] & ~in_2_V[40] & ~in_3_V[40] & ~weight_0_15_V_read[40]);
wire tmp_15_41;
assign tmp_15_41 = (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_15_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_15_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_15_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_15_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_15_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_15_V_read[41]) | (1 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_15_V_read[41]) | (0 &  in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_15_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_15_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_15_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_15_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_15_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_15_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_15_V_read[41]) | (1 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_15_V_read[41]) | (0 &  in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_15_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_15_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_15_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_15_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_15_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_15_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_15_V_read[41]) | (0 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_15_V_read[41]) | (1 & ~in_V[41] &  in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_15_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] &  weight_0_15_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] &  in_3_V[41] & ~weight_0_15_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] &  weight_0_15_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] &  in_2_V[41] & ~in_3_V[41] & ~weight_0_15_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] &  weight_0_15_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] &  in_3_V[41] & ~weight_0_15_V_read[41]) | (0 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] &  weight_0_15_V_read[41]) | (1 & ~in_V[41] & ~in_1_V[41] & ~in_2_V[41] & ~in_3_V[41] & ~weight_0_15_V_read[41]);
wire tmp_15_42;
assign tmp_15_42 = (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_15_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_15_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_15_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_15_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_15_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_15_V_read[42]) | (1 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_15_V_read[42]) | (0 &  in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_15_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_15_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_15_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_15_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_15_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_15_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_15_V_read[42]) | (1 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_15_V_read[42]) | (0 &  in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_15_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_15_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_15_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_15_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_15_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_15_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_15_V_read[42]) | (0 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_15_V_read[42]) | (1 & ~in_V[42] &  in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_15_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] &  weight_0_15_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] &  in_3_V[42] & ~weight_0_15_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] &  weight_0_15_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] &  in_2_V[42] & ~in_3_V[42] & ~weight_0_15_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] &  weight_0_15_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] &  in_3_V[42] & ~weight_0_15_V_read[42]) | (0 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] &  weight_0_15_V_read[42]) | (1 & ~in_V[42] & ~in_1_V[42] & ~in_2_V[42] & ~in_3_V[42] & ~weight_0_15_V_read[42]);
wire tmp_15_43;
assign tmp_15_43 = (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_15_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_15_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_15_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_15_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_15_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_15_V_read[43]) | (1 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_15_V_read[43]) | (0 &  in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_15_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_15_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_15_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_15_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_15_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_15_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_15_V_read[43]) | (1 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_15_V_read[43]) | (0 &  in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_15_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_15_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_15_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_15_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_15_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_15_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_15_V_read[43]) | (0 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_15_V_read[43]) | (1 & ~in_V[43] &  in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_15_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] &  weight_0_15_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] &  in_3_V[43] & ~weight_0_15_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] &  weight_0_15_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] &  in_2_V[43] & ~in_3_V[43] & ~weight_0_15_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] &  weight_0_15_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] &  in_3_V[43] & ~weight_0_15_V_read[43]) | (0 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] &  weight_0_15_V_read[43]) | (1 & ~in_V[43] & ~in_1_V[43] & ~in_2_V[43] & ~in_3_V[43] & ~weight_0_15_V_read[43]);
wire tmp_15_44;
assign tmp_15_44 = (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_15_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_15_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_15_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_15_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_15_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_15_V_read[44]) | (1 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_15_V_read[44]) | (0 &  in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_15_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_15_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_15_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_15_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_15_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_15_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_15_V_read[44]) | (1 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_15_V_read[44]) | (0 &  in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_15_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_15_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_15_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_15_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_15_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_15_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_15_V_read[44]) | (0 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_15_V_read[44]) | (1 & ~in_V[44] &  in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_15_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] &  weight_0_15_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] &  in_3_V[44] & ~weight_0_15_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] &  weight_0_15_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] &  in_2_V[44] & ~in_3_V[44] & ~weight_0_15_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] &  weight_0_15_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] &  in_3_V[44] & ~weight_0_15_V_read[44]) | (0 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] &  weight_0_15_V_read[44]) | (1 & ~in_V[44] & ~in_1_V[44] & ~in_2_V[44] & ~in_3_V[44] & ~weight_0_15_V_read[44]);
wire tmp_15_45;
assign tmp_15_45 = (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_15_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_15_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_15_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_15_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_15_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_15_V_read[45]) | (1 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_15_V_read[45]) | (0 &  in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_15_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_15_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_15_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_15_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_15_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_15_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_15_V_read[45]) | (1 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_15_V_read[45]) | (0 &  in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_15_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_15_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_15_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_15_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_15_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_15_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_15_V_read[45]) | (0 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_15_V_read[45]) | (1 & ~in_V[45] &  in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_15_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] &  weight_0_15_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] &  in_3_V[45] & ~weight_0_15_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] &  weight_0_15_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] &  in_2_V[45] & ~in_3_V[45] & ~weight_0_15_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] &  weight_0_15_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] &  in_3_V[45] & ~weight_0_15_V_read[45]) | (0 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] &  weight_0_15_V_read[45]) | (1 & ~in_V[45] & ~in_1_V[45] & ~in_2_V[45] & ~in_3_V[45] & ~weight_0_15_V_read[45]);
wire tmp_15_47;
assign tmp_15_47 = (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_15_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_15_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_15_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_15_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_15_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_15_V_read[47]) | (1 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_15_V_read[47]) | (0 &  in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_15_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_15_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_15_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_15_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_15_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_15_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_15_V_read[47]) | (1 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_15_V_read[47]) | (0 &  in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_15_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_15_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_15_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_15_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_15_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_15_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_15_V_read[47]) | (0 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_15_V_read[47]) | (1 & ~in_V[47] &  in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_15_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] &  weight_0_15_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] &  in_3_V[47] & ~weight_0_15_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] &  weight_0_15_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] &  in_2_V[47] & ~in_3_V[47] & ~weight_0_15_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] &  weight_0_15_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] &  in_3_V[47] & ~weight_0_15_V_read[47]) | (0 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] &  weight_0_15_V_read[47]) | (1 & ~in_V[47] & ~in_1_V[47] & ~in_2_V[47] & ~in_3_V[47] & ~weight_0_15_V_read[47]);
wire tmp_15_48;
assign tmp_15_48 = (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_15_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_15_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_15_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_15_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_15_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_15_V_read[48]) | (1 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_15_V_read[48]) | (0 &  in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_15_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_15_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_15_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_15_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_15_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_15_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_15_V_read[48]) | (1 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_15_V_read[48]) | (0 &  in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_15_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_15_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_15_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_15_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_15_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_15_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_15_V_read[48]) | (0 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_15_V_read[48]) | (1 & ~in_V[48] &  in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_15_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] &  weight_0_15_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] &  in_3_V[48] & ~weight_0_15_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] &  weight_0_15_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] &  in_2_V[48] & ~in_3_V[48] & ~weight_0_15_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] &  weight_0_15_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] &  in_3_V[48] & ~weight_0_15_V_read[48]) | (0 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] &  weight_0_15_V_read[48]) | (1 & ~in_V[48] & ~in_1_V[48] & ~in_2_V[48] & ~in_3_V[48] & ~weight_0_15_V_read[48]);
wire tmp_15_49;
assign tmp_15_49 = (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_15_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_15_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_15_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_15_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_15_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_15_V_read[49]) | (1 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_15_V_read[49]) | (0 &  in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_15_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_15_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_15_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_15_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_15_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_15_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_15_V_read[49]) | (1 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_15_V_read[49]) | (0 &  in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_15_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_15_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_15_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_15_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_15_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_15_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_15_V_read[49]) | (0 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_15_V_read[49]) | (1 & ~in_V[49] &  in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_15_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] &  weight_0_15_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] &  in_3_V[49] & ~weight_0_15_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] &  weight_0_15_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] &  in_2_V[49] & ~in_3_V[49] & ~weight_0_15_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] &  weight_0_15_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] &  in_3_V[49] & ~weight_0_15_V_read[49]) | (0 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] &  weight_0_15_V_read[49]) | (1 & ~in_V[49] & ~in_1_V[49] & ~in_2_V[49] & ~in_3_V[49] & ~weight_0_15_V_read[49]);
wire tmp_15_50;
assign tmp_15_50 = (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_15_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_15_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_15_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_15_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_15_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_15_V_read[50]) | (1 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_15_V_read[50]) | (0 &  in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_15_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_15_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_15_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_15_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_15_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_15_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_15_V_read[50]) | (1 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_15_V_read[50]) | (0 &  in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_15_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_15_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_15_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_15_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_15_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_15_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_15_V_read[50]) | (0 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_15_V_read[50]) | (1 & ~in_V[50] &  in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_15_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] &  weight_0_15_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] &  in_3_V[50] & ~weight_0_15_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] &  weight_0_15_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] &  in_2_V[50] & ~in_3_V[50] & ~weight_0_15_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] &  weight_0_15_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] &  in_3_V[50] & ~weight_0_15_V_read[50]) | (0 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] &  weight_0_15_V_read[50]) | (1 & ~in_V[50] & ~in_1_V[50] & ~in_2_V[50] & ~in_3_V[50] & ~weight_0_15_V_read[50]);
wire tmp_15_51;
assign tmp_15_51 = (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_15_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_15_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_15_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_15_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_15_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_15_V_read[51]) | (1 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_15_V_read[51]) | (0 &  in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_15_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_15_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_15_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_15_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_15_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_15_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_15_V_read[51]) | (1 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_15_V_read[51]) | (0 &  in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_15_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_15_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_15_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_15_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_15_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_15_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_15_V_read[51]) | (0 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_15_V_read[51]) | (1 & ~in_V[51] &  in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_15_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] &  weight_0_15_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] &  in_3_V[51] & ~weight_0_15_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] &  weight_0_15_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] &  in_2_V[51] & ~in_3_V[51] & ~weight_0_15_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] &  weight_0_15_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] &  in_3_V[51] & ~weight_0_15_V_read[51]) | (0 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] &  weight_0_15_V_read[51]) | (1 & ~in_V[51] & ~in_1_V[51] & ~in_2_V[51] & ~in_3_V[51] & ~weight_0_15_V_read[51]);
wire tmp_15_52;
assign tmp_15_52 = (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_15_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_15_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_15_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_15_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_15_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_15_V_read[52]) | (1 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_15_V_read[52]) | (0 &  in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_15_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_15_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_15_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_15_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_15_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_15_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_15_V_read[52]) | (1 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_15_V_read[52]) | (0 &  in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_15_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_15_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_15_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_15_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_15_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_15_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_15_V_read[52]) | (0 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_15_V_read[52]) | (1 & ~in_V[52] &  in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_15_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] &  weight_0_15_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] &  in_3_V[52] & ~weight_0_15_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] &  weight_0_15_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] &  in_2_V[52] & ~in_3_V[52] & ~weight_0_15_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] &  weight_0_15_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] &  in_3_V[52] & ~weight_0_15_V_read[52]) | (0 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] &  weight_0_15_V_read[52]) | (1 & ~in_V[52] & ~in_1_V[52] & ~in_2_V[52] & ~in_3_V[52] & ~weight_0_15_V_read[52]);
wire tmp_15_53;
assign tmp_15_53 = (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_15_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_15_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_15_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_15_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_15_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_15_V_read[53]) | (1 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_15_V_read[53]) | (0 &  in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_15_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_15_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_15_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_15_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_15_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_15_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_15_V_read[53]) | (1 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_15_V_read[53]) | (0 &  in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_15_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_15_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_15_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_15_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_15_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_15_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_15_V_read[53]) | (0 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_15_V_read[53]) | (1 & ~in_V[53] &  in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_15_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] &  weight_0_15_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] &  in_3_V[53] & ~weight_0_15_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] &  weight_0_15_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] &  in_2_V[53] & ~in_3_V[53] & ~weight_0_15_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] &  weight_0_15_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] &  in_3_V[53] & ~weight_0_15_V_read[53]) | (0 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] &  weight_0_15_V_read[53]) | (1 & ~in_V[53] & ~in_1_V[53] & ~in_2_V[53] & ~in_3_V[53] & ~weight_0_15_V_read[53]);
wire tmp_15_54;
assign tmp_15_54 = (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_15_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_15_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_15_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_15_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_15_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_15_V_read[54]) | (1 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_15_V_read[54]) | (0 &  in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_15_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_15_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_15_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_15_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_15_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_15_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_15_V_read[54]) | (1 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_15_V_read[54]) | (0 &  in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_15_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_15_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_15_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_15_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_15_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_15_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_15_V_read[54]) | (0 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_15_V_read[54]) | (1 & ~in_V[54] &  in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_15_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] &  weight_0_15_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] &  in_3_V[54] & ~weight_0_15_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] &  weight_0_15_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] &  in_2_V[54] & ~in_3_V[54] & ~weight_0_15_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] &  weight_0_15_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] &  in_3_V[54] & ~weight_0_15_V_read[54]) | (0 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] &  weight_0_15_V_read[54]) | (1 & ~in_V[54] & ~in_1_V[54] & ~in_2_V[54] & ~in_3_V[54] & ~weight_0_15_V_read[54]);
wire tmp_15_55;
assign tmp_15_55 = (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_15_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_15_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_15_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_15_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_15_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_15_V_read[55]) | (1 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_15_V_read[55]) | (0 &  in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_15_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_15_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_15_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_15_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_15_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_15_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_15_V_read[55]) | (1 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_15_V_read[55]) | (0 &  in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_15_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_15_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_15_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_15_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_15_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_15_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_15_V_read[55]) | (0 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_15_V_read[55]) | (1 & ~in_V[55] &  in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_15_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] &  weight_0_15_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] &  in_3_V[55] & ~weight_0_15_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] &  weight_0_15_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] &  in_2_V[55] & ~in_3_V[55] & ~weight_0_15_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] &  weight_0_15_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] &  in_3_V[55] & ~weight_0_15_V_read[55]) | (0 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] &  weight_0_15_V_read[55]) | (1 & ~in_V[55] & ~in_1_V[55] & ~in_2_V[55] & ~in_3_V[55] & ~weight_0_15_V_read[55]);
wire tmp_15_56;
assign tmp_15_56 = (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_15_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_15_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_15_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_15_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_15_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_15_V_read[56]) | (1 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_15_V_read[56]) | (0 &  in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_15_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_15_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_15_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_15_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_15_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_15_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_15_V_read[56]) | (1 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_15_V_read[56]) | (0 &  in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_15_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_15_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_15_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_15_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_15_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_15_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_15_V_read[56]) | (0 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_15_V_read[56]) | (1 & ~in_V[56] &  in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_15_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] &  weight_0_15_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] &  in_3_V[56] & ~weight_0_15_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] &  weight_0_15_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] &  in_2_V[56] & ~in_3_V[56] & ~weight_0_15_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] &  weight_0_15_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] &  in_3_V[56] & ~weight_0_15_V_read[56]) | (0 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] &  weight_0_15_V_read[56]) | (1 & ~in_V[56] & ~in_1_V[56] & ~in_2_V[56] & ~in_3_V[56] & ~weight_0_15_V_read[56]);
wire tmp_15_57;
assign tmp_15_57 = (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_15_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_15_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_15_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_15_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_15_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_15_V_read[57]) | (1 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_15_V_read[57]) | (0 &  in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_15_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_15_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_15_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_15_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_15_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_15_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_15_V_read[57]) | (1 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_15_V_read[57]) | (0 &  in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_15_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_15_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_15_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_15_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_15_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_15_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_15_V_read[57]) | (0 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_15_V_read[57]) | (1 & ~in_V[57] &  in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_15_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] &  weight_0_15_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] &  in_3_V[57] & ~weight_0_15_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] &  weight_0_15_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] &  in_2_V[57] & ~in_3_V[57] & ~weight_0_15_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] &  weight_0_15_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] &  in_3_V[57] & ~weight_0_15_V_read[57]) | (0 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] &  weight_0_15_V_read[57]) | (1 & ~in_V[57] & ~in_1_V[57] & ~in_2_V[57] & ~in_3_V[57] & ~weight_0_15_V_read[57]);
wire tmp_15_58;
assign tmp_15_58 = (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_15_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_15_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_15_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_15_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_15_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_15_V_read[58]) | (1 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_15_V_read[58]) | (0 &  in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_15_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_15_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_15_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_15_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_15_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_15_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_15_V_read[58]) | (1 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_15_V_read[58]) | (0 &  in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_15_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_15_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_15_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_15_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_15_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_15_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_15_V_read[58]) | (0 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_15_V_read[58]) | (1 & ~in_V[58] &  in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_15_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] &  weight_0_15_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] &  in_3_V[58] & ~weight_0_15_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] &  weight_0_15_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] &  in_2_V[58] & ~in_3_V[58] & ~weight_0_15_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] &  weight_0_15_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] &  in_3_V[58] & ~weight_0_15_V_read[58]) | (0 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] &  weight_0_15_V_read[58]) | (1 & ~in_V[58] & ~in_1_V[58] & ~in_2_V[58] & ~in_3_V[58] & ~weight_0_15_V_read[58]);
wire tmp_15_59;
assign tmp_15_59 = (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_15_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_15_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_15_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_15_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_15_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_15_V_read[59]) | (1 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_15_V_read[59]) | (0 &  in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_15_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_15_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_15_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_15_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_15_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_15_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_15_V_read[59]) | (1 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_15_V_read[59]) | (0 &  in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_15_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_15_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_15_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_15_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_15_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_15_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_15_V_read[59]) | (0 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_15_V_read[59]) | (1 & ~in_V[59] &  in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_15_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] &  weight_0_15_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] &  in_3_V[59] & ~weight_0_15_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] &  weight_0_15_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] &  in_2_V[59] & ~in_3_V[59] & ~weight_0_15_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] &  weight_0_15_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] &  in_3_V[59] & ~weight_0_15_V_read[59]) | (0 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] &  weight_0_15_V_read[59]) | (1 & ~in_V[59] & ~in_1_V[59] & ~in_2_V[59] & ~in_3_V[59] & ~weight_0_15_V_read[59]);
wire tmp_15_60;
assign tmp_15_60 = (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_15_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_15_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_15_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_15_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_15_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_15_V_read[60]) | (1 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_15_V_read[60]) | (0 &  in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_15_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_15_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_15_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_15_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_15_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_15_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_15_V_read[60]) | (1 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_15_V_read[60]) | (0 &  in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_15_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_15_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_15_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_15_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_15_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_15_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_15_V_read[60]) | (0 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_15_V_read[60]) | (1 & ~in_V[60] &  in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_15_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] &  weight_0_15_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] &  in_3_V[60] & ~weight_0_15_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] &  weight_0_15_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] &  in_2_V[60] & ~in_3_V[60] & ~weight_0_15_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] &  weight_0_15_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] &  in_3_V[60] & ~weight_0_15_V_read[60]) | (0 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] &  weight_0_15_V_read[60]) | (1 & ~in_V[60] & ~in_1_V[60] & ~in_2_V[60] & ~in_3_V[60] & ~weight_0_15_V_read[60]);
wire tmp_15_62;
assign tmp_15_62 = (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_15_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_15_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_15_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_15_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_15_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_15_V_read[62]) | (1 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_15_V_read[62]) | (0 &  in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_15_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_15_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_15_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_15_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_15_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_15_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_15_V_read[62]) | (1 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_15_V_read[62]) | (0 &  in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_15_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_15_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_15_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_15_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_15_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_15_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_15_V_read[62]) | (0 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_15_V_read[62]) | (1 & ~in_V[62] &  in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_15_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] &  weight_0_15_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] &  in_3_V[62] & ~weight_0_15_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] &  weight_0_15_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] &  in_2_V[62] & ~in_3_V[62] & ~weight_0_15_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] &  weight_0_15_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] &  in_3_V[62] & ~weight_0_15_V_read[62]) | (0 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] &  weight_0_15_V_read[62]) | (1 & ~in_V[62] & ~in_1_V[62] & ~in_2_V[62] & ~in_3_V[62] & ~weight_0_15_V_read[62]);
wire tmp_15_63;
assign tmp_15_63 = (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_15_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_15_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_15_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_15_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_15_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_15_V_read[63]) | (1 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_15_V_read[63]) | (0 &  in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_15_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_15_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_15_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_15_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_15_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_15_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_15_V_read[63]) | (1 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_15_V_read[63]) | (0 &  in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_15_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_15_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_15_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_15_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_15_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_15_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_15_V_read[63]) | (0 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_15_V_read[63]) | (1 & ~in_V[63] &  in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_15_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] &  weight_0_15_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] &  in_3_V[63] & ~weight_0_15_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] &  weight_0_15_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] &  in_2_V[63] & ~in_3_V[63] & ~weight_0_15_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] &  weight_0_15_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] &  in_3_V[63] & ~weight_0_15_V_read[63]) | (0 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] &  weight_0_15_V_read[63]) | (1 & ~in_V[63] & ~in_1_V[63] & ~in_2_V[63] & ~in_3_V[63] & ~weight_0_15_V_read[63]);
wire tmp_15_64;
assign tmp_15_64 = (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_15_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_15_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_15_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_15_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_15_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_15_V_read[64]) | (1 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_15_V_read[64]) | (0 &  in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_15_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_15_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_15_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_15_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_15_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_15_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_15_V_read[64]) | (1 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_15_V_read[64]) | (0 &  in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_15_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_15_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_15_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_15_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_15_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_15_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_15_V_read[64]) | (0 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_15_V_read[64]) | (1 & ~in_V[64] &  in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_15_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] &  weight_0_15_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] &  in_3_V[64] & ~weight_0_15_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] &  weight_0_15_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] &  in_2_V[64] & ~in_3_V[64] & ~weight_0_15_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] &  weight_0_15_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] &  in_3_V[64] & ~weight_0_15_V_read[64]) | (0 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] &  weight_0_15_V_read[64]) | (1 & ~in_V[64] & ~in_1_V[64] & ~in_2_V[64] & ~in_3_V[64] & ~weight_0_15_V_read[64]);
wire tmp_15_65;
assign tmp_15_65 = (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_15_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_15_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_15_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_15_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_15_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_15_V_read[65]) | (1 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_15_V_read[65]) | (0 &  in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_15_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_15_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_15_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_15_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_15_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_15_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_15_V_read[65]) | (1 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_15_V_read[65]) | (0 &  in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_15_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_15_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_15_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_15_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_15_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_15_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_15_V_read[65]) | (0 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_15_V_read[65]) | (1 & ~in_V[65] &  in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_15_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] &  weight_0_15_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] &  in_3_V[65] & ~weight_0_15_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] &  weight_0_15_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] &  in_2_V[65] & ~in_3_V[65] & ~weight_0_15_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] &  weight_0_15_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] &  in_3_V[65] & ~weight_0_15_V_read[65]) | (0 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] &  weight_0_15_V_read[65]) | (1 & ~in_V[65] & ~in_1_V[65] & ~in_2_V[65] & ~in_3_V[65] & ~weight_0_15_V_read[65]);
wire tmp_15_66;
assign tmp_15_66 = (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_15_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_15_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_15_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_15_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_15_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_15_V_read[66]) | (1 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_15_V_read[66]) | (0 &  in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_15_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_15_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_15_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_15_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_15_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_15_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_15_V_read[66]) | (1 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_15_V_read[66]) | (0 &  in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_15_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_15_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_15_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_15_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_15_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_15_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_15_V_read[66]) | (0 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_15_V_read[66]) | (1 & ~in_V[66] &  in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_15_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] &  weight_0_15_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] &  in_3_V[66] & ~weight_0_15_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] &  weight_0_15_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] &  in_2_V[66] & ~in_3_V[66] & ~weight_0_15_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] &  weight_0_15_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] &  in_3_V[66] & ~weight_0_15_V_read[66]) | (0 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] &  weight_0_15_V_read[66]) | (1 & ~in_V[66] & ~in_1_V[66] & ~in_2_V[66] & ~in_3_V[66] & ~weight_0_15_V_read[66]);
wire tmp_15_67;
assign tmp_15_67 = (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_15_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_15_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_15_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_15_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_15_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_15_V_read[67]) | (1 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_15_V_read[67]) | (0 &  in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_15_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_15_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_15_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_15_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_15_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_15_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_15_V_read[67]) | (1 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_15_V_read[67]) | (0 &  in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_15_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_15_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_15_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_15_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_15_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_15_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_15_V_read[67]) | (0 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_15_V_read[67]) | (1 & ~in_V[67] &  in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_15_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] &  weight_0_15_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] &  in_3_V[67] & ~weight_0_15_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] &  weight_0_15_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] &  in_2_V[67] & ~in_3_V[67] & ~weight_0_15_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] &  weight_0_15_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] &  in_3_V[67] & ~weight_0_15_V_read[67]) | (0 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] &  weight_0_15_V_read[67]) | (1 & ~in_V[67] & ~in_1_V[67] & ~in_2_V[67] & ~in_3_V[67] & ~weight_0_15_V_read[67]);
wire tmp_15_68;
assign tmp_15_68 = (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_15_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_15_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_15_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_15_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_15_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_15_V_read[68]) | (1 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_15_V_read[68]) | (0 &  in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_15_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_15_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_15_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_15_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_15_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_15_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_15_V_read[68]) | (1 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_15_V_read[68]) | (0 &  in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_15_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_15_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_15_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_15_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_15_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_15_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_15_V_read[68]) | (0 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_15_V_read[68]) | (1 & ~in_V[68] &  in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_15_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] &  weight_0_15_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] &  in_3_V[68] & ~weight_0_15_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] &  weight_0_15_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] &  in_2_V[68] & ~in_3_V[68] & ~weight_0_15_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] &  weight_0_15_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] &  in_3_V[68] & ~weight_0_15_V_read[68]) | (0 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] &  weight_0_15_V_read[68]) | (1 & ~in_V[68] & ~in_1_V[68] & ~in_2_V[68] & ~in_3_V[68] & ~weight_0_15_V_read[68]);
wire tmp_15_69;
assign tmp_15_69 = (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_15_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_15_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_15_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_15_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_15_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_15_V_read[69]) | (1 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_15_V_read[69]) | (0 &  in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_15_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_15_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_15_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_15_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_15_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_15_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_15_V_read[69]) | (1 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_15_V_read[69]) | (0 &  in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_15_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_15_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_15_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_15_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_15_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_15_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_15_V_read[69]) | (0 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_15_V_read[69]) | (1 & ~in_V[69] &  in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_15_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] &  weight_0_15_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] &  in_3_V[69] & ~weight_0_15_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] &  weight_0_15_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] &  in_2_V[69] & ~in_3_V[69] & ~weight_0_15_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] &  weight_0_15_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] &  in_3_V[69] & ~weight_0_15_V_read[69]) | (0 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] &  weight_0_15_V_read[69]) | (1 & ~in_V[69] & ~in_1_V[69] & ~in_2_V[69] & ~in_3_V[69] & ~weight_0_15_V_read[69]);
wire tmp_15_70;
assign tmp_15_70 = (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_15_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_15_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_15_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_15_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_15_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_15_V_read[70]) | (1 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_15_V_read[70]) | (0 &  in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_15_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_15_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_15_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_15_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_15_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_15_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_15_V_read[70]) | (1 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_15_V_read[70]) | (0 &  in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_15_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_15_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_15_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_15_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_15_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_15_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_15_V_read[70]) | (0 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_15_V_read[70]) | (1 & ~in_V[70] &  in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_15_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] &  weight_0_15_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] &  in_3_V[70] & ~weight_0_15_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] &  weight_0_15_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] &  in_2_V[70] & ~in_3_V[70] & ~weight_0_15_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] &  weight_0_15_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] &  in_3_V[70] & ~weight_0_15_V_read[70]) | (0 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] &  weight_0_15_V_read[70]) | (1 & ~in_V[70] & ~in_1_V[70] & ~in_2_V[70] & ~in_3_V[70] & ~weight_0_15_V_read[70]);
assign ap_return_15 = {tmp_15_0,tmp_15_1,tmp_15_2,tmp_15_3,tmp_15_4,tmp_15_5,tmp_15_6,tmp_15_7,tmp_15_8,tmp_15_9,tmp_15_10,1'b0,tmp_15_12,tmp_15_13,tmp_15_14,tmp_15_15,tmp_15_16,tmp_15_17,tmp_15_18,tmp_15_19,tmp_15_20,tmp_15_21,tmp_15_22,tmp_15_23,tmp_15_24,tmp_15_25,tmp_15_26,tmp_15_27,tmp_15_28,tmp_15_29,tmp_15_30,1'b0,1'b0,tmp_15_33,1'b0,tmp_15_35,1'b0,tmp_15_37,tmp_15_38,tmp_15_39,tmp_15_40,tmp_15_41,tmp_15_42,tmp_15_43,tmp_15_44,tmp_15_45,1'b0,tmp_15_47,tmp_15_48,tmp_15_49,tmp_15_50,tmp_15_51,tmp_15_52,tmp_15_53,tmp_15_54,tmp_15_55,tmp_15_56,tmp_15_57,tmp_15_58,tmp_15_59,tmp_15_60,1'b0,tmp_15_62,tmp_15_63,tmp_15_64,tmp_15_65,tmp_15_66,tmp_15_67,tmp_15_68,tmp_15_69,tmp_15_70,1'b0};
endmodule